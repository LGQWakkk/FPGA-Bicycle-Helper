`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/06/07 22:46:39
// Design Name: 
// Module Name: map_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//注意：这里面输入的坐标以地图为原点
//为了节约带宽资源
//map_x需要除以8
//map_y由于范围在0-239所以使用8位来表示
//最终大小是14位

module map_rom(
    input wire clk,
	input wire [13:0] addr,//map_y[7:0]  map_x[8:3]  {8,6}
	output reg [7:0] data  //输出的一行像素
    );
	
	reg [13:0] addr_reg;
	
	always@(posedge clk)begin
		addr_reg<=addr;
	end
	
	always@(*)begin
		case(addr_reg)
14'h0000:data=8'hFF;
14'h0001:data=8'hFF;
14'h0002:data=8'hFF;
14'h0003:data=8'hC0;
14'h0004:data=8'h00;
14'h0005:data=8'h00;
14'h0006:data=8'h00;
14'h0007:data=8'h00;
14'h0008:data=8'h00;
14'h0009:data=8'h00;
14'h000a:data=8'h00;
14'h000b:data=8'h00;
14'h000c:data=8'h00;
14'h000d:data=8'h00;
14'h000e:data=8'h00;
14'h000f:data=8'h00;
14'h0010:data=8'h00;
14'h0011:data=8'h00;
14'h0012:data=8'h00;
14'h0013:data=8'h00;
14'h0014:data=8'h00;
14'h0015:data=8'h00;
14'h0016:data=8'h00;
14'h0017:data=8'h00;
14'h0018:data=8'h00;
14'h0019:data=8'h07;
14'h001a:data=8'hFF;
14'h001b:data=8'hFF;
14'h001c:data=8'hFF;
14'h001d:data=8'hFF;
14'h001e:data=8'hFF;
14'h001f:data=8'hFF;
14'h0020:data=8'hFF;
14'h0021:data=8'hFF;
14'h0022:data=8'hFF;
14'h0023:data=8'hFF;
14'h0024:data=8'hFF;
14'h0025:data=8'hFC;
14'h0026:data=8'h00;
14'h0027:data=8'h00;
14'h0040:data=8'hFF;
14'h0041:data=8'hFF;
14'h0042:data=8'hFF;
14'h0043:data=8'hC0;
14'h0044:data=8'h00;
14'h0045:data=8'h00;
14'h0046:data=8'h00;
14'h0047:data=8'h00;
14'h0048:data=8'h00;
14'h0049:data=8'h00;
14'h004a:data=8'h00;
14'h004b:data=8'h00;
14'h004c:data=8'h00;
14'h004d:data=8'h00;
14'h004e:data=8'h00;
14'h004f:data=8'h00;
14'h0050:data=8'h00;
14'h0051:data=8'h00;
14'h0052:data=8'h00;
14'h0053:data=8'h00;
14'h0054:data=8'h00;
14'h0055:data=8'h00;
14'h0056:data=8'h00;
14'h0057:data=8'h00;
14'h0058:data=8'h00;
14'h0059:data=8'h07;
14'h005a:data=8'hFF;
14'h005b:data=8'hFF;
14'h005c:data=8'hFF;
14'h005d:data=8'hFF;
14'h005e:data=8'hFF;
14'h005f:data=8'hFF;
14'h0060:data=8'hFF;
14'h0061:data=8'hFF;
14'h0062:data=8'hFF;
14'h0063:data=8'hFF;
14'h0064:data=8'hFF;
14'h0065:data=8'hFC;
14'h0066:data=8'h00;
14'h0067:data=8'h00;
14'h0080:data=8'hFF;
14'h0081:data=8'hFF;
14'h0082:data=8'hFF;
14'h0083:data=8'hC0;
14'h0084:data=8'h00;
14'h0085:data=8'h00;
14'h0086:data=8'h00;
14'h0087:data=8'h00;
14'h0088:data=8'h00;
14'h0089:data=8'h00;
14'h008a:data=8'h00;
14'h008b:data=8'h00;
14'h008c:data=8'h00;
14'h008d:data=8'h00;
14'h008e:data=8'h00;
14'h008f:data=8'h00;
14'h0090:data=8'h00;
14'h0091:data=8'h00;
14'h0092:data=8'h00;
14'h0093:data=8'h00;
14'h0094:data=8'h00;
14'h0095:data=8'h00;
14'h0096:data=8'h00;
14'h0097:data=8'h00;
14'h0098:data=8'h00;
14'h0099:data=8'h07;
14'h009a:data=8'hFF;
14'h009b:data=8'hFF;
14'h009c:data=8'hFF;
14'h009d:data=8'hFF;
14'h009e:data=8'hFF;
14'h009f:data=8'hFF;
14'h00a0:data=8'hFF;
14'h00a1:data=8'hFF;
14'h00a2:data=8'hFF;
14'h00a3:data=8'hFF;
14'h00a4:data=8'hFF;
14'h00a5:data=8'hFC;
14'h00a6:data=8'h00;
14'h00a7:data=8'h00;
14'h00c0:data=8'hFF;
14'h00c1:data=8'hFF;
14'h00c2:data=8'hFF;
14'h00c3:data=8'hC0;
14'h00c4:data=8'h00;
14'h00c5:data=8'h00;
14'h00c6:data=8'h00;
14'h00c7:data=8'h00;
14'h00c8:data=8'h00;
14'h00c9:data=8'h00;
14'h00ca:data=8'h00;
14'h00cb:data=8'h00;
14'h00cc:data=8'h00;
14'h00cd:data=8'h00;
14'h00ce:data=8'h00;
14'h00cf:data=8'h00;
14'h00d0:data=8'h00;
14'h00d1:data=8'h00;
14'h00d2:data=8'h00;
14'h00d3:data=8'h00;
14'h00d4:data=8'h00;
14'h00d5:data=8'h00;
14'h00d6:data=8'h00;
14'h00d7:data=8'h00;
14'h00d8:data=8'h00;
14'h00d9:data=8'h07;
14'h00da:data=8'hFF;
14'h00db:data=8'hFF;
14'h00dc:data=8'hFF;
14'h00dd:data=8'hFF;
14'h00de:data=8'hFF;
14'h00df:data=8'hFF;
14'h00e0:data=8'hFF;
14'h00e1:data=8'hFF;
14'h00e2:data=8'hFF;
14'h00e3:data=8'hFF;
14'h00e4:data=8'hFF;
14'h00e5:data=8'hFC;
14'h00e6:data=8'h00;
14'h00e7:data=8'h00;
14'h0100:data=8'hFF;
14'h0101:data=8'hFF;
14'h0102:data=8'hFF;
14'h0103:data=8'hC0;
14'h0104:data=8'h00;
14'h0105:data=8'h00;
14'h0106:data=8'h00;
14'h0107:data=8'h00;
14'h0108:data=8'h00;
14'h0109:data=8'h00;
14'h010a:data=8'h00;
14'h010b:data=8'h00;
14'h010c:data=8'h00;
14'h010d:data=8'h00;
14'h010e:data=8'h00;
14'h010f:data=8'h00;
14'h0110:data=8'h00;
14'h0111:data=8'h00;
14'h0112:data=8'h00;
14'h0113:data=8'h00;
14'h0114:data=8'h00;
14'h0115:data=8'h00;
14'h0116:data=8'h00;
14'h0117:data=8'h00;
14'h0118:data=8'h00;
14'h0119:data=8'h07;
14'h011a:data=8'hFF;
14'h011b:data=8'hFF;
14'h011c:data=8'hFF;
14'h011d:data=8'hFF;
14'h011e:data=8'hFF;
14'h011f:data=8'hFF;
14'h0120:data=8'hFF;
14'h0121:data=8'hFF;
14'h0122:data=8'hFF;
14'h0123:data=8'hFF;
14'h0124:data=8'hFF;
14'h0125:data=8'hFC;
14'h0126:data=8'h00;
14'h0127:data=8'h00;
14'h0140:data=8'hFF;
14'h0141:data=8'hFF;
14'h0142:data=8'hFF;
14'h0143:data=8'hC0;
14'h0144:data=8'h00;
14'h0145:data=8'h00;
14'h0146:data=8'h00;
14'h0147:data=8'h00;
14'h0148:data=8'h00;
14'h0149:data=8'h00;
14'h014a:data=8'h00;
14'h014b:data=8'h00;
14'h014c:data=8'h00;
14'h014d:data=8'h00;
14'h014e:data=8'h00;
14'h014f:data=8'h00;
14'h0150:data=8'h00;
14'h0151:data=8'h00;
14'h0152:data=8'h00;
14'h0153:data=8'h00;
14'h0154:data=8'h00;
14'h0155:data=8'h00;
14'h0156:data=8'h00;
14'h0157:data=8'h00;
14'h0158:data=8'h00;
14'h0159:data=8'h07;
14'h015a:data=8'hFF;
14'h015b:data=8'hFF;
14'h015c:data=8'hFF;
14'h015d:data=8'hFF;
14'h015e:data=8'hFF;
14'h015f:data=8'hFF;
14'h0160:data=8'hFF;
14'h0161:data=8'hFF;
14'h0162:data=8'hFF;
14'h0163:data=8'hFF;
14'h0164:data=8'hFF;
14'h0165:data=8'hFC;
14'h0166:data=8'h00;
14'h0167:data=8'h00;
14'h0180:data=8'hFF;
14'h0181:data=8'hFF;
14'h0182:data=8'hFF;
14'h0183:data=8'hC0;
14'h0184:data=8'h00;
14'h0185:data=8'h00;
14'h0186:data=8'h00;
14'h0187:data=8'h00;
14'h0188:data=8'h00;
14'h0189:data=8'h00;
14'h018a:data=8'h00;
14'h018b:data=8'h00;
14'h018c:data=8'h00;
14'h018d:data=8'h00;
14'h018e:data=8'h00;
14'h018f:data=8'h00;
14'h0190:data=8'h00;
14'h0191:data=8'h00;
14'h0192:data=8'h00;
14'h0193:data=8'h00;
14'h0194:data=8'h00;
14'h0195:data=8'h00;
14'h0196:data=8'h00;
14'h0197:data=8'h00;
14'h0198:data=8'h00;
14'h0199:data=8'h07;
14'h019a:data=8'hFF;
14'h019b:data=8'hFF;
14'h019c:data=8'hFF;
14'h019d:data=8'hFF;
14'h019e:data=8'hFF;
14'h019f:data=8'hFF;
14'h01a0:data=8'hFF;
14'h01a1:data=8'hFF;
14'h01a2:data=8'hFF;
14'h01a3:data=8'hFF;
14'h01a4:data=8'hFF;
14'h01a5:data=8'hFC;
14'h01a6:data=8'h00;
14'h01a7:data=8'h00;
14'h01c0:data=8'h01;
14'h01c1:data=8'hFF;
14'h01c2:data=8'hFF;
14'h01c3:data=8'hC0;
14'h01c4:data=8'h00;
14'h01c5:data=8'h00;
14'h01c6:data=8'h00;
14'h01c7:data=8'h00;
14'h01c8:data=8'h00;
14'h01c9:data=8'h00;
14'h01ca:data=8'h00;
14'h01cb:data=8'h00;
14'h01cc:data=8'h00;
14'h01cd:data=8'h00;
14'h01ce:data=8'h00;
14'h01cf:data=8'h00;
14'h01d0:data=8'h00;
14'h01d1:data=8'h00;
14'h01d2:data=8'h00;
14'h01d3:data=8'h00;
14'h01d4:data=8'h00;
14'h01d5:data=8'h00;
14'h01d6:data=8'h00;
14'h01d7:data=8'h00;
14'h01d8:data=8'h00;
14'h01d9:data=8'h07;
14'h01da:data=8'hFF;
14'h01db:data=8'hFF;
14'h01dc:data=8'hFC;
14'h01dd:data=8'h00;
14'h01de:data=8'h00;
14'h01df:data=8'h00;
14'h01e0:data=8'h00;
14'h01e1:data=8'h00;
14'h01e2:data=8'h1F;
14'h01e3:data=8'hFF;
14'h01e4:data=8'hFF;
14'h01e5:data=8'hFC;
14'h01e6:data=8'h00;
14'h01e7:data=8'h00;
14'h0200:data=8'h01;
14'h0201:data=8'hFF;
14'h0202:data=8'hFF;
14'h0203:data=8'hC0;
14'h0204:data=8'h00;
14'h0205:data=8'h00;
14'h0206:data=8'h00;
14'h0207:data=8'h00;
14'h0208:data=8'h00;
14'h0209:data=8'h00;
14'h020a:data=8'h00;
14'h020b:data=8'h00;
14'h020c:data=8'h00;
14'h020d:data=8'h00;
14'h020e:data=8'h00;
14'h020f:data=8'h00;
14'h0210:data=8'h00;
14'h0211:data=8'h00;
14'h0212:data=8'h00;
14'h0213:data=8'h00;
14'h0214:data=8'h00;
14'h0215:data=8'h00;
14'h0216:data=8'h00;
14'h0217:data=8'h00;
14'h0218:data=8'h00;
14'h0219:data=8'h07;
14'h021a:data=8'hFF;
14'h021b:data=8'hFF;
14'h021c:data=8'hFC;
14'h021d:data=8'h00;
14'h021e:data=8'h00;
14'h021f:data=8'h00;
14'h0220:data=8'h00;
14'h0221:data=8'h00;
14'h0222:data=8'h1F;
14'h0223:data=8'hFF;
14'h0224:data=8'hFF;
14'h0225:data=8'hFC;
14'h0226:data=8'h00;
14'h0227:data=8'h00;
14'h0240:data=8'h01;
14'h0241:data=8'hFF;
14'h0242:data=8'hFF;
14'h0243:data=8'hC0;
14'h0244:data=8'h00;
14'h0245:data=8'h00;
14'h0246:data=8'h00;
14'h0247:data=8'h00;
14'h0248:data=8'h00;
14'h0249:data=8'h00;
14'h024a:data=8'h00;
14'h024b:data=8'h00;
14'h024c:data=8'h00;
14'h024d:data=8'h00;
14'h024e:data=8'h00;
14'h024f:data=8'h00;
14'h0250:data=8'h00;
14'h0251:data=8'h00;
14'h0252:data=8'h00;
14'h0253:data=8'h00;
14'h0254:data=8'h00;
14'h0255:data=8'h00;
14'h0256:data=8'h00;
14'h0257:data=8'h00;
14'h0258:data=8'h00;
14'h0259:data=8'h07;
14'h025a:data=8'hFF;
14'h025b:data=8'hFF;
14'h025c:data=8'hFC;
14'h025d:data=8'h00;
14'h025e:data=8'h00;
14'h025f:data=8'h00;
14'h0260:data=8'h00;
14'h0261:data=8'h00;
14'h0262:data=8'h1F;
14'h0263:data=8'hFF;
14'h0264:data=8'hFF;
14'h0265:data=8'hFC;
14'h0266:data=8'h00;
14'h0267:data=8'h00;
14'h0280:data=8'h01;
14'h0281:data=8'hFF;
14'h0282:data=8'hFF;
14'h0283:data=8'hC0;
14'h0284:data=8'h00;
14'h0285:data=8'h00;
14'h0286:data=8'h00;
14'h0287:data=8'h00;
14'h0288:data=8'h00;
14'h0289:data=8'h00;
14'h028a:data=8'h00;
14'h028b:data=8'h00;
14'h028c:data=8'h00;
14'h028d:data=8'h00;
14'h028e:data=8'h00;
14'h028f:data=8'h00;
14'h0290:data=8'h00;
14'h0291:data=8'h00;
14'h0292:data=8'h00;
14'h0293:data=8'h00;
14'h0294:data=8'h00;
14'h0295:data=8'h00;
14'h0296:data=8'h00;
14'h0297:data=8'h00;
14'h0298:data=8'h00;
14'h0299:data=8'h07;
14'h029a:data=8'hFF;
14'h029b:data=8'hFF;
14'h029c:data=8'hFC;
14'h029d:data=8'h00;
14'h029e:data=8'h00;
14'h029f:data=8'h00;
14'h02a0:data=8'h00;
14'h02a1:data=8'h00;
14'h02a2:data=8'h1F;
14'h02a3:data=8'hFF;
14'h02a4:data=8'hFF;
14'h02a5:data=8'hFC;
14'h02a6:data=8'h00;
14'h02a7:data=8'h00;
14'h02c0:data=8'h01;
14'h02c1:data=8'hFF;
14'h02c2:data=8'hFF;
14'h02c3:data=8'hC0;
14'h02c4:data=8'h00;
14'h02c5:data=8'h00;
14'h02c6:data=8'h00;
14'h02c7:data=8'h00;
14'h02c8:data=8'h00;
14'h02c9:data=8'h00;
14'h02ca:data=8'h00;
14'h02cb:data=8'h00;
14'h02cc:data=8'h00;
14'h02cd:data=8'h00;
14'h02ce:data=8'h00;
14'h02cf:data=8'h00;
14'h02d0:data=8'h00;
14'h02d1:data=8'h00;
14'h02d2:data=8'h00;
14'h02d3:data=8'h00;
14'h02d4:data=8'h00;
14'h02d5:data=8'h00;
14'h02d6:data=8'h00;
14'h02d7:data=8'h00;
14'h02d8:data=8'h00;
14'h02d9:data=8'h07;
14'h02da:data=8'hFF;
14'h02db:data=8'hFF;
14'h02dc:data=8'hFC;
14'h02dd:data=8'h00;
14'h02de:data=8'h00;
14'h02df:data=8'h00;
14'h02e0:data=8'h00;
14'h02e1:data=8'h00;
14'h02e2:data=8'h1F;
14'h02e3:data=8'hFF;
14'h02e4:data=8'hFF;
14'h02e5:data=8'hFC;
14'h02e6:data=8'h00;
14'h02e7:data=8'h00;
14'h0300:data=8'h01;
14'h0301:data=8'hFF;
14'h0302:data=8'hFF;
14'h0303:data=8'hC0;
14'h0304:data=8'h00;
14'h0305:data=8'h00;
14'h0306:data=8'h00;
14'h0307:data=8'h00;
14'h0308:data=8'h00;
14'h0309:data=8'h00;
14'h030a:data=8'h00;
14'h030b:data=8'h00;
14'h030c:data=8'h00;
14'h030d:data=8'h00;
14'h030e:data=8'h00;
14'h030f:data=8'h00;
14'h0310:data=8'h00;
14'h0311:data=8'h00;
14'h0312:data=8'h00;
14'h0313:data=8'h00;
14'h0314:data=8'h00;
14'h0315:data=8'h00;
14'h0316:data=8'h00;
14'h0317:data=8'h00;
14'h0318:data=8'h00;
14'h0319:data=8'h07;
14'h031a:data=8'hFF;
14'h031b:data=8'hFF;
14'h031c:data=8'hFC;
14'h031d:data=8'h00;
14'h031e:data=8'h00;
14'h031f:data=8'h00;
14'h0320:data=8'h00;
14'h0321:data=8'h00;
14'h0322:data=8'h1F;
14'h0323:data=8'hFF;
14'h0324:data=8'hFF;
14'h0325:data=8'hFC;
14'h0326:data=8'h00;
14'h0327:data=8'h00;
14'h0340:data=8'h01;
14'h0341:data=8'hFF;
14'h0342:data=8'hFF;
14'h0343:data=8'hC0;
14'h0344:data=8'h00;
14'h0345:data=8'h00;
14'h0346:data=8'h00;
14'h0347:data=8'h00;
14'h0348:data=8'h00;
14'h0349:data=8'h00;
14'h034a:data=8'h00;
14'h034b:data=8'h00;
14'h034c:data=8'h00;
14'h034d:data=8'h00;
14'h034e:data=8'h00;
14'h034f:data=8'h00;
14'h0350:data=8'h00;
14'h0351:data=8'h00;
14'h0352:data=8'h00;
14'h0353:data=8'h00;
14'h0354:data=8'h00;
14'h0355:data=8'h00;
14'h0356:data=8'h00;
14'h0357:data=8'h00;
14'h0358:data=8'h00;
14'h0359:data=8'h07;
14'h035a:data=8'hFF;
14'h035b:data=8'hFF;
14'h035c:data=8'hFC;
14'h035d:data=8'h00;
14'h035e:data=8'h00;
14'h035f:data=8'h00;
14'h0360:data=8'h00;
14'h0361:data=8'h00;
14'h0362:data=8'h1F;
14'h0363:data=8'hFF;
14'h0364:data=8'hFF;
14'h0365:data=8'hFC;
14'h0366:data=8'h00;
14'h0367:data=8'h00;
14'h0380:data=8'h01;
14'h0381:data=8'hFF;
14'h0382:data=8'hFF;
14'h0383:data=8'hC0;
14'h0384:data=8'h00;
14'h0385:data=8'h00;
14'h0386:data=8'h00;
14'h0387:data=8'h00;
14'h0388:data=8'h00;
14'h0389:data=8'h00;
14'h038a:data=8'h00;
14'h038b:data=8'h00;
14'h038c:data=8'h00;
14'h038d:data=8'h00;
14'h038e:data=8'h00;
14'h038f:data=8'h00;
14'h0390:data=8'h00;
14'h0391:data=8'h00;
14'h0392:data=8'h00;
14'h0393:data=8'h00;
14'h0394:data=8'h00;
14'h0395:data=8'h00;
14'h0396:data=8'h00;
14'h0397:data=8'h00;
14'h0398:data=8'h00;
14'h0399:data=8'h07;
14'h039a:data=8'hFF;
14'h039b:data=8'hFF;
14'h039c:data=8'hFC;
14'h039d:data=8'h00;
14'h039e:data=8'h00;
14'h039f:data=8'h00;
14'h03a0:data=8'h00;
14'h03a1:data=8'h00;
14'h03a2:data=8'h1F;
14'h03a3:data=8'hFF;
14'h03a4:data=8'hFF;
14'h03a5:data=8'hFC;
14'h03a6:data=8'h00;
14'h03a7:data=8'h00;
14'h03c0:data=8'h01;
14'h03c1:data=8'hFF;
14'h03c2:data=8'hFF;
14'h03c3:data=8'hC0;
14'h03c4:data=8'h00;
14'h03c5:data=8'h00;
14'h03c6:data=8'h00;
14'h03c7:data=8'h00;
14'h03c8:data=8'h00;
14'h03c9:data=8'h00;
14'h03ca:data=8'h00;
14'h03cb:data=8'h00;
14'h03cc:data=8'h00;
14'h03cd:data=8'h00;
14'h03ce:data=8'h00;
14'h03cf:data=8'h00;
14'h03d0:data=8'h00;
14'h03d1:data=8'h00;
14'h03d2:data=8'h00;
14'h03d3:data=8'h00;
14'h03d4:data=8'h00;
14'h03d5:data=8'h00;
14'h03d6:data=8'h00;
14'h03d7:data=8'h00;
14'h03d8:data=8'h00;
14'h03d9:data=8'h07;
14'h03da:data=8'hFF;
14'h03db:data=8'hFF;
14'h03dc:data=8'hFC;
14'h03dd:data=8'h00;
14'h03de:data=8'h00;
14'h03df:data=8'h00;
14'h03e0:data=8'h00;
14'h03e1:data=8'h00;
14'h03e2:data=8'h1F;
14'h03e3:data=8'hFF;
14'h03e4:data=8'hFF;
14'h03e5:data=8'hFC;
14'h03e6:data=8'h00;
14'h03e7:data=8'h00;
14'h0400:data=8'h01;
14'h0401:data=8'hFF;
14'h0402:data=8'hFF;
14'h0403:data=8'hC0;
14'h0404:data=8'h00;
14'h0405:data=8'h00;
14'h0406:data=8'h00;
14'h0407:data=8'h00;
14'h0408:data=8'h00;
14'h0409:data=8'h00;
14'h040a:data=8'h00;
14'h040b:data=8'h00;
14'h040c:data=8'h00;
14'h040d:data=8'h00;
14'h040e:data=8'h00;
14'h040f:data=8'h00;
14'h0410:data=8'h00;
14'h0411:data=8'h00;
14'h0412:data=8'h00;
14'h0413:data=8'h00;
14'h0414:data=8'h00;
14'h0415:data=8'h00;
14'h0416:data=8'h00;
14'h0417:data=8'h00;
14'h0418:data=8'h00;
14'h0419:data=8'h07;
14'h041a:data=8'hFF;
14'h041b:data=8'hFF;
14'h041c:data=8'hFC;
14'h041d:data=8'h00;
14'h041e:data=8'h00;
14'h041f:data=8'h00;
14'h0420:data=8'h00;
14'h0421:data=8'h00;
14'h0422:data=8'h1F;
14'h0423:data=8'hFF;
14'h0424:data=8'hFF;
14'h0425:data=8'hFC;
14'h0426:data=8'h00;
14'h0427:data=8'h00;
14'h0440:data=8'h01;
14'h0441:data=8'hFF;
14'h0442:data=8'hFF;
14'h0443:data=8'hC0;
14'h0444:data=8'h00;
14'h0445:data=8'h00;
14'h0446:data=8'h00;
14'h0447:data=8'h00;
14'h0448:data=8'h00;
14'h0449:data=8'h00;
14'h044a:data=8'h00;
14'h044b:data=8'h00;
14'h044c:data=8'h00;
14'h044d:data=8'h00;
14'h044e:data=8'h00;
14'h044f:data=8'h00;
14'h0450:data=8'h00;
14'h0451:data=8'h00;
14'h0452:data=8'h00;
14'h0453:data=8'h00;
14'h0454:data=8'h00;
14'h0455:data=8'h00;
14'h0456:data=8'h00;
14'h0457:data=8'h00;
14'h0458:data=8'h00;
14'h0459:data=8'h07;
14'h045a:data=8'hFF;
14'h045b:data=8'hFF;
14'h045c:data=8'hFC;
14'h045d:data=8'h00;
14'h045e:data=8'h00;
14'h045f:data=8'h00;
14'h0460:data=8'h00;
14'h0461:data=8'h00;
14'h0462:data=8'h1F;
14'h0463:data=8'hFF;
14'h0464:data=8'hFF;
14'h0465:data=8'hFC;
14'h0466:data=8'h00;
14'h0467:data=8'h00;
14'h0480:data=8'h01;
14'h0481:data=8'hFF;
14'h0482:data=8'hFF;
14'h0483:data=8'hC0;
14'h0484:data=8'h00;
14'h0485:data=8'h00;
14'h0486:data=8'h00;
14'h0487:data=8'h00;
14'h0488:data=8'h00;
14'h0489:data=8'h00;
14'h048a:data=8'h00;
14'h048b:data=8'h00;
14'h048c:data=8'h00;
14'h048d:data=8'h00;
14'h048e:data=8'h00;
14'h048f:data=8'h00;
14'h0490:data=8'h00;
14'h0491:data=8'h00;
14'h0492:data=8'h00;
14'h0493:data=8'h00;
14'h0494:data=8'h00;
14'h0495:data=8'h00;
14'h0496:data=8'h00;
14'h0497:data=8'h00;
14'h0498:data=8'h00;
14'h0499:data=8'h07;
14'h049a:data=8'hFF;
14'h049b:data=8'hFF;
14'h049c:data=8'hFC;
14'h049d:data=8'h00;
14'h049e:data=8'h00;
14'h049f:data=8'h00;
14'h04a0:data=8'h00;
14'h04a1:data=8'h00;
14'h04a2:data=8'h1F;
14'h04a3:data=8'hFF;
14'h04a4:data=8'hFF;
14'h04a5:data=8'hFC;
14'h04a6:data=8'h00;
14'h04a7:data=8'h00;
14'h04c0:data=8'h01;
14'h04c1:data=8'hFF;
14'h04c2:data=8'hFF;
14'h04c3:data=8'hC0;
14'h04c4:data=8'h00;
14'h04c5:data=8'h00;
14'h04c6:data=8'h00;
14'h04c7:data=8'h00;
14'h04c8:data=8'h00;
14'h04c9:data=8'h00;
14'h04ca:data=8'h00;
14'h04cb:data=8'h00;
14'h04cc:data=8'h00;
14'h04cd:data=8'h00;
14'h04ce:data=8'h00;
14'h04cf:data=8'h00;
14'h04d0:data=8'h00;
14'h04d1:data=8'h00;
14'h04d2:data=8'h00;
14'h04d3:data=8'h00;
14'h04d4:data=8'h00;
14'h04d5:data=8'h00;
14'h04d6:data=8'h00;
14'h04d7:data=8'h00;
14'h04d8:data=8'h00;
14'h04d9:data=8'h07;
14'h04da:data=8'hFF;
14'h04db:data=8'hFF;
14'h04dc:data=8'hFC;
14'h04dd:data=8'h00;
14'h04de:data=8'h00;
14'h04df:data=8'h00;
14'h04e0:data=8'h00;
14'h04e1:data=8'h00;
14'h04e2:data=8'h1F;
14'h04e3:data=8'hFF;
14'h04e4:data=8'hFF;
14'h04e5:data=8'hFC;
14'h04e6:data=8'h00;
14'h04e7:data=8'h00;
14'h0500:data=8'h01;
14'h0501:data=8'hFF;
14'h0502:data=8'hFF;
14'h0503:data=8'hC0;
14'h0504:data=8'h00;
14'h0505:data=8'h00;
14'h0506:data=8'h00;
14'h0507:data=8'h00;
14'h0508:data=8'h00;
14'h0509:data=8'h00;
14'h050a:data=8'h00;
14'h050b:data=8'h00;
14'h050c:data=8'h00;
14'h050d:data=8'h00;
14'h050e:data=8'h00;
14'h050f:data=8'h00;
14'h0510:data=8'h00;
14'h0511:data=8'h00;
14'h0512:data=8'h00;
14'h0513:data=8'h00;
14'h0514:data=8'h00;
14'h0515:data=8'h00;
14'h0516:data=8'h00;
14'h0517:data=8'h00;
14'h0518:data=8'h00;
14'h0519:data=8'h07;
14'h051a:data=8'hFF;
14'h051b:data=8'hFF;
14'h051c:data=8'hFC;
14'h051d:data=8'h00;
14'h051e:data=8'h00;
14'h051f:data=8'h00;
14'h0520:data=8'h00;
14'h0521:data=8'h00;
14'h0522:data=8'h1F;
14'h0523:data=8'hFF;
14'h0524:data=8'hFF;
14'h0525:data=8'hFC;
14'h0526:data=8'h00;
14'h0527:data=8'h00;
14'h0540:data=8'h01;
14'h0541:data=8'hFF;
14'h0542:data=8'hFF;
14'h0543:data=8'hC0;
14'h0544:data=8'h00;
14'h0545:data=8'h00;
14'h0546:data=8'h00;
14'h0547:data=8'h00;
14'h0548:data=8'h00;
14'h0549:data=8'h00;
14'h054a:data=8'h00;
14'h054b:data=8'h00;
14'h054c:data=8'h00;
14'h054d:data=8'h00;
14'h054e:data=8'h00;
14'h054f:data=8'h00;
14'h0550:data=8'h00;
14'h0551:data=8'h00;
14'h0552:data=8'h00;
14'h0553:data=8'h00;
14'h0554:data=8'h00;
14'h0555:data=8'h00;
14'h0556:data=8'h00;
14'h0557:data=8'h00;
14'h0558:data=8'h00;
14'h0559:data=8'h07;
14'h055a:data=8'hFF;
14'h055b:data=8'hFF;
14'h055c:data=8'hFC;
14'h055d:data=8'h00;
14'h055e:data=8'h00;
14'h055f:data=8'h00;
14'h0560:data=8'h00;
14'h0561:data=8'h00;
14'h0562:data=8'h1F;
14'h0563:data=8'hFF;
14'h0564:data=8'hFF;
14'h0565:data=8'hFC;
14'h0566:data=8'h00;
14'h0567:data=8'h00;
14'h0580:data=8'h01;
14'h0581:data=8'hFF;
14'h0582:data=8'hFF;
14'h0583:data=8'hC0;
14'h0584:data=8'h00;
14'h0585:data=8'h00;
14'h0586:data=8'h00;
14'h0587:data=8'h00;
14'h0588:data=8'h00;
14'h0589:data=8'h00;
14'h058a:data=8'h00;
14'h058b:data=8'h00;
14'h058c:data=8'h00;
14'h058d:data=8'h00;
14'h058e:data=8'h00;
14'h058f:data=8'h00;
14'h0590:data=8'h00;
14'h0591:data=8'h00;
14'h0592:data=8'h00;
14'h0593:data=8'h00;
14'h0594:data=8'h00;
14'h0595:data=8'h00;
14'h0596:data=8'h00;
14'h0597:data=8'h00;
14'h0598:data=8'h00;
14'h0599:data=8'h07;
14'h059a:data=8'hFF;
14'h059b:data=8'hFF;
14'h059c:data=8'hFC;
14'h059d:data=8'h00;
14'h059e:data=8'h00;
14'h059f:data=8'h00;
14'h05a0:data=8'h00;
14'h05a1:data=8'h00;
14'h05a2:data=8'h1F;
14'h05a3:data=8'hFF;
14'h05a4:data=8'hFF;
14'h05a5:data=8'hFC;
14'h05a6:data=8'h00;
14'h05a7:data=8'h00;
14'h05c0:data=8'h01;
14'h05c1:data=8'hFF;
14'h05c2:data=8'hFF;
14'h05c3:data=8'hC0;
14'h05c4:data=8'h00;
14'h05c5:data=8'h00;
14'h05c6:data=8'h00;
14'h05c7:data=8'h00;
14'h05c8:data=8'h00;
14'h05c9:data=8'h00;
14'h05ca:data=8'h00;
14'h05cb:data=8'h00;
14'h05cc:data=8'h00;
14'h05cd:data=8'h00;
14'h05ce:data=8'h00;
14'h05cf:data=8'h00;
14'h05d0:data=8'h00;
14'h05d1:data=8'h00;
14'h05d2:data=8'h00;
14'h05d3:data=8'h00;
14'h05d4:data=8'h00;
14'h05d5:data=8'h00;
14'h05d6:data=8'h00;
14'h05d7:data=8'h00;
14'h05d8:data=8'h00;
14'h05d9:data=8'h07;
14'h05da:data=8'hFF;
14'h05db:data=8'hFF;
14'h05dc:data=8'hFC;
14'h05dd:data=8'h00;
14'h05de:data=8'h00;
14'h05df:data=8'h00;
14'h05e0:data=8'h00;
14'h05e1:data=8'h00;
14'h05e2:data=8'h1F;
14'h05e3:data=8'hFF;
14'h05e4:data=8'hFF;
14'h05e5:data=8'hFC;
14'h05e6:data=8'h00;
14'h05e7:data=8'h00;
14'h0600:data=8'h01;
14'h0601:data=8'hFF;
14'h0602:data=8'hFF;
14'h0603:data=8'hC0;
14'h0604:data=8'h00;
14'h0605:data=8'h00;
14'h0606:data=8'h00;
14'h0607:data=8'h00;
14'h0608:data=8'h00;
14'h0609:data=8'h00;
14'h060a:data=8'h00;
14'h060b:data=8'h00;
14'h060c:data=8'h00;
14'h060d:data=8'h00;
14'h060e:data=8'h00;
14'h060f:data=8'h00;
14'h0610:data=8'h00;
14'h0611:data=8'h00;
14'h0612:data=8'h00;
14'h0613:data=8'h00;
14'h0614:data=8'h00;
14'h0615:data=8'h00;
14'h0616:data=8'h00;
14'h0617:data=8'h00;
14'h0618:data=8'h00;
14'h0619:data=8'h07;
14'h061a:data=8'hFF;
14'h061b:data=8'hFF;
14'h061c:data=8'hFC;
14'h061d:data=8'h00;
14'h061e:data=8'h00;
14'h061f:data=8'h00;
14'h0620:data=8'h00;
14'h0621:data=8'h00;
14'h0622:data=8'h1F;
14'h0623:data=8'hFF;
14'h0624:data=8'hFF;
14'h0625:data=8'hFC;
14'h0626:data=8'h00;
14'h0627:data=8'h00;
14'h0640:data=8'h01;
14'h0641:data=8'hFF;
14'h0642:data=8'hFF;
14'h0643:data=8'hC0;
14'h0644:data=8'h00;
14'h0645:data=8'h00;
14'h0646:data=8'h00;
14'h0647:data=8'h00;
14'h0648:data=8'h00;
14'h0649:data=8'h00;
14'h064a:data=8'h00;
14'h064b:data=8'h00;
14'h064c:data=8'h00;
14'h064d:data=8'h00;
14'h064e:data=8'h00;
14'h064f:data=8'h00;
14'h0650:data=8'h00;
14'h0651:data=8'h00;
14'h0652:data=8'h00;
14'h0653:data=8'h00;
14'h0654:data=8'h00;
14'h0655:data=8'h00;
14'h0656:data=8'h00;
14'h0657:data=8'h00;
14'h0658:data=8'h00;
14'h0659:data=8'h07;
14'h065a:data=8'hFF;
14'h065b:data=8'hFF;
14'h065c:data=8'hFC;
14'h065d:data=8'h00;
14'h065e:data=8'h00;
14'h065f:data=8'h00;
14'h0660:data=8'h00;
14'h0661:data=8'h00;
14'h0662:data=8'h1F;
14'h0663:data=8'hFF;
14'h0664:data=8'hFF;
14'h0665:data=8'hFC;
14'h0666:data=8'h00;
14'h0667:data=8'h00;
14'h0680:data=8'h01;
14'h0681:data=8'hFF;
14'h0682:data=8'hFF;
14'h0683:data=8'hC0;
14'h0684:data=8'h00;
14'h0685:data=8'h00;
14'h0686:data=8'h00;
14'h0687:data=8'h00;
14'h0688:data=8'h00;
14'h0689:data=8'h00;
14'h068a:data=8'h00;
14'h068b:data=8'h00;
14'h068c:data=8'h00;
14'h068d:data=8'h00;
14'h068e:data=8'h00;
14'h068f:data=8'h00;
14'h0690:data=8'h00;
14'h0691:data=8'h00;
14'h0692:data=8'h00;
14'h0693:data=8'h00;
14'h0694:data=8'h00;
14'h0695:data=8'h00;
14'h0696:data=8'h00;
14'h0697:data=8'h00;
14'h0698:data=8'h00;
14'h0699:data=8'h07;
14'h069a:data=8'hFF;
14'h069b:data=8'hFF;
14'h069c:data=8'hFC;
14'h069d:data=8'h00;
14'h069e:data=8'h00;
14'h069f:data=8'h00;
14'h06a0:data=8'h00;
14'h06a1:data=8'h00;
14'h06a2:data=8'h1F;
14'h06a3:data=8'hFF;
14'h06a4:data=8'hFF;
14'h06a5:data=8'hFC;
14'h06a6:data=8'h00;
14'h06a7:data=8'h00;
14'h06c0:data=8'h01;
14'h06c1:data=8'hFF;
14'h06c2:data=8'hFF;
14'h06c3:data=8'hC0;
14'h06c4:data=8'h00;
14'h06c5:data=8'h00;
14'h06c6:data=8'h00;
14'h06c7:data=8'h00;
14'h06c8:data=8'h00;
14'h06c9:data=8'h00;
14'h06ca:data=8'h00;
14'h06cb:data=8'h00;
14'h06cc:data=8'h00;
14'h06cd:data=8'h00;
14'h06ce:data=8'h00;
14'h06cf:data=8'h00;
14'h06d0:data=8'h00;
14'h06d1:data=8'h00;
14'h06d2:data=8'h00;
14'h06d3:data=8'h00;
14'h06d4:data=8'h00;
14'h06d5:data=8'h00;
14'h06d6:data=8'h00;
14'h06d7:data=8'h00;
14'h06d8:data=8'h00;
14'h06d9:data=8'h07;
14'h06da:data=8'hFF;
14'h06db:data=8'hFF;
14'h06dc:data=8'hFC;
14'h06dd:data=8'h00;
14'h06de:data=8'h00;
14'h06df:data=8'h00;
14'h06e0:data=8'h00;
14'h06e1:data=8'h00;
14'h06e2:data=8'h1F;
14'h06e3:data=8'hFF;
14'h06e4:data=8'hFF;
14'h06e5:data=8'hFC;
14'h06e6:data=8'h00;
14'h06e7:data=8'h00;
14'h0700:data=8'h01;
14'h0701:data=8'hFF;
14'h0702:data=8'hFF;
14'h0703:data=8'hC0;
14'h0704:data=8'h00;
14'h0705:data=8'h00;
14'h0706:data=8'h00;
14'h0707:data=8'h00;
14'h0708:data=8'h00;
14'h0709:data=8'h00;
14'h070a:data=8'h00;
14'h070b:data=8'h00;
14'h070c:data=8'h00;
14'h070d:data=8'h00;
14'h070e:data=8'h00;
14'h070f:data=8'h00;
14'h0710:data=8'h00;
14'h0711:data=8'h00;
14'h0712:data=8'h00;
14'h0713:data=8'h00;
14'h0714:data=8'h00;
14'h0715:data=8'h00;
14'h0716:data=8'h00;
14'h0717:data=8'h00;
14'h0718:data=8'h00;
14'h0719:data=8'h07;
14'h071a:data=8'hFF;
14'h071b:data=8'hFF;
14'h071c:data=8'hFC;
14'h071d:data=8'h00;
14'h071e:data=8'h00;
14'h071f:data=8'h00;
14'h0720:data=8'h00;
14'h0721:data=8'h00;
14'h0722:data=8'h1F;
14'h0723:data=8'hFF;
14'h0724:data=8'hFF;
14'h0725:data=8'hFC;
14'h0726:data=8'h00;
14'h0727:data=8'h00;
14'h0740:data=8'h01;
14'h0741:data=8'hFF;
14'h0742:data=8'hFF;
14'h0743:data=8'hC0;
14'h0744:data=8'h00;
14'h0745:data=8'h00;
14'h0746:data=8'h00;
14'h0747:data=8'h00;
14'h0748:data=8'h00;
14'h0749:data=8'h00;
14'h074a:data=8'h00;
14'h074b:data=8'h00;
14'h074c:data=8'h00;
14'h074d:data=8'h00;
14'h074e:data=8'h00;
14'h074f:data=8'h00;
14'h0750:data=8'h00;
14'h0751:data=8'h00;
14'h0752:data=8'h00;
14'h0753:data=8'h00;
14'h0754:data=8'h00;
14'h0755:data=8'h00;
14'h0756:data=8'h00;
14'h0757:data=8'h00;
14'h0758:data=8'h00;
14'h0759:data=8'h07;
14'h075a:data=8'hFF;
14'h075b:data=8'hFF;
14'h075c:data=8'hFC;
14'h075d:data=8'h00;
14'h075e:data=8'h00;
14'h075f:data=8'h00;
14'h0760:data=8'h00;
14'h0761:data=8'h00;
14'h0762:data=8'h1F;
14'h0763:data=8'hFF;
14'h0764:data=8'hFF;
14'h0765:data=8'hFC;
14'h0766:data=8'h00;
14'h0767:data=8'h00;
14'h0780:data=8'h01;
14'h0781:data=8'hFF;
14'h0782:data=8'hFF;
14'h0783:data=8'hC0;
14'h0784:data=8'h00;
14'h0785:data=8'h00;
14'h0786:data=8'h00;
14'h0787:data=8'h00;
14'h0788:data=8'h00;
14'h0789:data=8'h00;
14'h078a:data=8'h00;
14'h078b:data=8'h00;
14'h078c:data=8'h00;
14'h078d:data=8'h00;
14'h078e:data=8'h00;
14'h078f:data=8'h00;
14'h0790:data=8'h00;
14'h0791:data=8'h00;
14'h0792:data=8'h00;
14'h0793:data=8'h00;
14'h0794:data=8'h00;
14'h0795:data=8'h00;
14'h0796:data=8'h00;
14'h0797:data=8'h00;
14'h0798:data=8'h00;
14'h0799:data=8'h07;
14'h079a:data=8'hFF;
14'h079b:data=8'hFF;
14'h079c:data=8'hFC;
14'h079d:data=8'h00;
14'h079e:data=8'h00;
14'h079f:data=8'h00;
14'h07a0:data=8'h00;
14'h07a1:data=8'h00;
14'h07a2:data=8'h1F;
14'h07a3:data=8'hFF;
14'h07a4:data=8'hFF;
14'h07a5:data=8'hFC;
14'h07a6:data=8'h00;
14'h07a7:data=8'h00;
14'h07c0:data=8'h01;
14'h07c1:data=8'hFF;
14'h07c2:data=8'hFF;
14'h07c3:data=8'hC0;
14'h07c4:data=8'h00;
14'h07c5:data=8'h00;
14'h07c6:data=8'h00;
14'h07c7:data=8'h00;
14'h07c8:data=8'h00;
14'h07c9:data=8'h00;
14'h07ca:data=8'h00;
14'h07cb:data=8'h00;
14'h07cc:data=8'h00;
14'h07cd:data=8'h00;
14'h07ce:data=8'h00;
14'h07cf:data=8'h00;
14'h07d0:data=8'h00;
14'h07d1:data=8'h00;
14'h07d2:data=8'h00;
14'h07d3:data=8'h00;
14'h07d4:data=8'h00;
14'h07d5:data=8'h00;
14'h07d6:data=8'h00;
14'h07d7:data=8'h00;
14'h07d8:data=8'h00;
14'h07d9:data=8'h07;
14'h07da:data=8'hFF;
14'h07db:data=8'hFF;
14'h07dc:data=8'hFC;
14'h07dd:data=8'h00;
14'h07de:data=8'h00;
14'h07df:data=8'h00;
14'h07e0:data=8'h00;
14'h07e1:data=8'h00;
14'h07e2:data=8'h1F;
14'h07e3:data=8'hFF;
14'h07e4:data=8'hFF;
14'h07e5:data=8'hFC;
14'h07e6:data=8'h00;
14'h07e7:data=8'h00;
14'h0800:data=8'h01;
14'h0801:data=8'hFF;
14'h0802:data=8'hFF;
14'h0803:data=8'hC0;
14'h0804:data=8'h00;
14'h0805:data=8'h00;
14'h0806:data=8'h00;
14'h0807:data=8'h00;
14'h0808:data=8'h00;
14'h0809:data=8'h00;
14'h080a:data=8'h00;
14'h080b:data=8'h00;
14'h080c:data=8'h00;
14'h080d:data=8'h00;
14'h080e:data=8'h00;
14'h080f:data=8'h00;
14'h0810:data=8'h00;
14'h0811:data=8'h00;
14'h0812:data=8'h00;
14'h0813:data=8'h00;
14'h0814:data=8'h00;
14'h0815:data=8'h00;
14'h0816:data=8'h00;
14'h0817:data=8'h00;
14'h0818:data=8'h00;
14'h0819:data=8'h07;
14'h081a:data=8'hFF;
14'h081b:data=8'hFF;
14'h081c:data=8'hFC;
14'h081d:data=8'h00;
14'h081e:data=8'h00;
14'h081f:data=8'h00;
14'h0820:data=8'h00;
14'h0821:data=8'h00;
14'h0822:data=8'h1F;
14'h0823:data=8'hFF;
14'h0824:data=8'hFF;
14'h0825:data=8'hFC;
14'h0826:data=8'h00;
14'h0827:data=8'h00;
14'h0840:data=8'h01;
14'h0841:data=8'hFF;
14'h0842:data=8'hFF;
14'h0843:data=8'hC0;
14'h0844:data=8'h00;
14'h0845:data=8'h00;
14'h0846:data=8'h00;
14'h0847:data=8'h00;
14'h0848:data=8'h00;
14'h0849:data=8'h00;
14'h084a:data=8'h00;
14'h084b:data=8'h00;
14'h084c:data=8'h00;
14'h084d:data=8'h00;
14'h084e:data=8'h00;
14'h084f:data=8'h00;
14'h0850:data=8'h00;
14'h0851:data=8'h00;
14'h0852:data=8'h00;
14'h0853:data=8'h00;
14'h0854:data=8'h00;
14'h0855:data=8'h00;
14'h0856:data=8'h00;
14'h0857:data=8'h00;
14'h0858:data=8'h00;
14'h0859:data=8'h07;
14'h085a:data=8'hFF;
14'h085b:data=8'hFF;
14'h085c:data=8'hFC;
14'h085d:data=8'h00;
14'h085e:data=8'h00;
14'h085f:data=8'h00;
14'h0860:data=8'h00;
14'h0861:data=8'h00;
14'h0862:data=8'h1F;
14'h0863:data=8'hFF;
14'h0864:data=8'hFF;
14'h0865:data=8'hFC;
14'h0866:data=8'h00;
14'h0867:data=8'h00;
14'h0880:data=8'h01;
14'h0881:data=8'hFF;
14'h0882:data=8'hFF;
14'h0883:data=8'hC0;
14'h0884:data=8'h00;
14'h0885:data=8'h00;
14'h0886:data=8'h00;
14'h0887:data=8'h00;
14'h0888:data=8'h00;
14'h0889:data=8'h00;
14'h088a:data=8'h00;
14'h088b:data=8'h00;
14'h088c:data=8'h00;
14'h088d:data=8'h00;
14'h088e:data=8'h00;
14'h088f:data=8'h00;
14'h0890:data=8'h00;
14'h0891:data=8'h00;
14'h0892:data=8'h00;
14'h0893:data=8'h00;
14'h0894:data=8'h00;
14'h0895:data=8'h00;
14'h0896:data=8'h00;
14'h0897:data=8'h00;
14'h0898:data=8'h00;
14'h0899:data=8'h07;
14'h089a:data=8'hFF;
14'h089b:data=8'hFF;
14'h089c:data=8'hFC;
14'h089d:data=8'h00;
14'h089e:data=8'h00;
14'h089f:data=8'h00;
14'h08a0:data=8'h00;
14'h08a1:data=8'h00;
14'h08a2:data=8'h1F;
14'h08a3:data=8'hFF;
14'h08a4:data=8'hFF;
14'h08a5:data=8'hFC;
14'h08a6:data=8'h00;
14'h08a7:data=8'h00;
14'h08c0:data=8'h01;
14'h08c1:data=8'hFF;
14'h08c2:data=8'hFF;
14'h08c3:data=8'hC0;
14'h08c4:data=8'h00;
14'h08c5:data=8'h00;
14'h08c6:data=8'h00;
14'h08c7:data=8'h00;
14'h08c8:data=8'h00;
14'h08c9:data=8'h00;
14'h08ca:data=8'h00;
14'h08cb:data=8'h00;
14'h08cc:data=8'h00;
14'h08cd:data=8'h00;
14'h08ce:data=8'h00;
14'h08cf:data=8'h00;
14'h08d0:data=8'h00;
14'h08d1:data=8'h00;
14'h08d2:data=8'h00;
14'h08d3:data=8'h00;
14'h08d4:data=8'h00;
14'h08d5:data=8'h00;
14'h08d6:data=8'h00;
14'h08d7:data=8'h00;
14'h08d8:data=8'h00;
14'h08d9:data=8'h07;
14'h08da:data=8'hFF;
14'h08db:data=8'hFF;
14'h08dc:data=8'hFC;
14'h08dd:data=8'h00;
14'h08de:data=8'h00;
14'h08df:data=8'h00;
14'h08e0:data=8'h00;
14'h08e1:data=8'h00;
14'h08e2:data=8'h1F;
14'h08e3:data=8'hFF;
14'h08e4:data=8'hFF;
14'h08e5:data=8'hFC;
14'h08e6:data=8'h00;
14'h08e7:data=8'h00;
14'h0900:data=8'h01;
14'h0901:data=8'hFF;
14'h0902:data=8'hFF;
14'h0903:data=8'hC0;
14'h0904:data=8'h00;
14'h0905:data=8'h00;
14'h0906:data=8'h00;
14'h0907:data=8'h00;
14'h0908:data=8'h00;
14'h0909:data=8'h00;
14'h090a:data=8'h00;
14'h090b:data=8'h00;
14'h090c:data=8'h00;
14'h090d:data=8'h00;
14'h090e:data=8'h00;
14'h090f:data=8'h00;
14'h0910:data=8'h00;
14'h0911:data=8'h00;
14'h0912:data=8'h00;
14'h0913:data=8'h00;
14'h0914:data=8'h00;
14'h0915:data=8'h00;
14'h0916:data=8'h00;
14'h0917:data=8'h00;
14'h0918:data=8'h00;
14'h0919:data=8'h07;
14'h091a:data=8'hFF;
14'h091b:data=8'hFF;
14'h091c:data=8'hFC;
14'h091d:data=8'h00;
14'h091e:data=8'h00;
14'h091f:data=8'h00;
14'h0920:data=8'h00;
14'h0921:data=8'h00;
14'h0922:data=8'h1F;
14'h0923:data=8'hFF;
14'h0924:data=8'hFF;
14'h0925:data=8'hFC;
14'h0926:data=8'h00;
14'h0927:data=8'h00;
14'h0940:data=8'h01;
14'h0941:data=8'hFF;
14'h0942:data=8'hFF;
14'h0943:data=8'hC0;
14'h0944:data=8'h00;
14'h0945:data=8'h00;
14'h0946:data=8'h00;
14'h0947:data=8'h00;
14'h0948:data=8'h00;
14'h0949:data=8'h00;
14'h094a:data=8'h00;
14'h094b:data=8'h00;
14'h094c:data=8'h00;
14'h094d:data=8'h00;
14'h094e:data=8'h00;
14'h094f:data=8'h00;
14'h0950:data=8'h00;
14'h0951:data=8'h00;
14'h0952:data=8'h00;
14'h0953:data=8'h00;
14'h0954:data=8'h00;
14'h0955:data=8'h00;
14'h0956:data=8'h00;
14'h0957:data=8'h00;
14'h0958:data=8'h00;
14'h0959:data=8'h07;
14'h095a:data=8'hFF;
14'h095b:data=8'hFF;
14'h095c:data=8'hFC;
14'h095d:data=8'h00;
14'h095e:data=8'h00;
14'h095f:data=8'h00;
14'h0960:data=8'h00;
14'h0961:data=8'h00;
14'h0962:data=8'h1F;
14'h0963:data=8'hFF;
14'h0964:data=8'hFF;
14'h0965:data=8'hFC;
14'h0966:data=8'h00;
14'h0967:data=8'h00;
14'h0980:data=8'h01;
14'h0981:data=8'hFF;
14'h0982:data=8'hFF;
14'h0983:data=8'hC0;
14'h0984:data=8'h00;
14'h0985:data=8'h00;
14'h0986:data=8'h00;
14'h0987:data=8'h00;
14'h0988:data=8'h00;
14'h0989:data=8'h00;
14'h098a:data=8'h00;
14'h098b:data=8'h00;
14'h098c:data=8'h00;
14'h098d:data=8'h00;
14'h098e:data=8'h00;
14'h098f:data=8'h00;
14'h0990:data=8'h00;
14'h0991:data=8'h00;
14'h0992:data=8'h00;
14'h0993:data=8'h00;
14'h0994:data=8'h00;
14'h0995:data=8'h00;
14'h0996:data=8'h00;
14'h0997:data=8'h00;
14'h0998:data=8'h00;
14'h0999:data=8'h07;
14'h099a:data=8'hFF;
14'h099b:data=8'hFF;
14'h099c:data=8'hFC;
14'h099d:data=8'h00;
14'h099e:data=8'h00;
14'h099f:data=8'h00;
14'h09a0:data=8'h00;
14'h09a1:data=8'h00;
14'h09a2:data=8'h1F;
14'h09a3:data=8'hFF;
14'h09a4:data=8'hFF;
14'h09a5:data=8'hFC;
14'h09a6:data=8'h00;
14'h09a7:data=8'h00;
14'h09c0:data=8'h01;
14'h09c1:data=8'hFF;
14'h09c2:data=8'hFF;
14'h09c3:data=8'hC0;
14'h09c4:data=8'h00;
14'h09c5:data=8'h00;
14'h09c6:data=8'h00;
14'h09c7:data=8'h00;
14'h09c8:data=8'h00;
14'h09c9:data=8'h00;
14'h09ca:data=8'h00;
14'h09cb:data=8'h00;
14'h09cc:data=8'h00;
14'h09cd:data=8'h00;
14'h09ce:data=8'h00;
14'h09cf:data=8'h00;
14'h09d0:data=8'h00;
14'h09d1:data=8'h00;
14'h09d2:data=8'h00;
14'h09d3:data=8'h00;
14'h09d4:data=8'h00;
14'h09d5:data=8'h00;
14'h09d6:data=8'h00;
14'h09d7:data=8'h00;
14'h09d8:data=8'h00;
14'h09d9:data=8'h07;
14'h09da:data=8'hFF;
14'h09db:data=8'hFF;
14'h09dc:data=8'hFC;
14'h09dd:data=8'h00;
14'h09de:data=8'h00;
14'h09df:data=8'h00;
14'h09e0:data=8'h00;
14'h09e1:data=8'h00;
14'h09e2:data=8'h1F;
14'h09e3:data=8'hFF;
14'h09e4:data=8'hFF;
14'h09e5:data=8'hFC;
14'h09e6:data=8'h00;
14'h09e7:data=8'h00;
14'h0a00:data=8'h01;
14'h0a01:data=8'hFF;
14'h0a02:data=8'hFF;
14'h0a03:data=8'hC0;
14'h0a04:data=8'h00;
14'h0a05:data=8'h00;
14'h0a06:data=8'h00;
14'h0a07:data=8'h00;
14'h0a08:data=8'h00;
14'h0a09:data=8'h00;
14'h0a0a:data=8'h00;
14'h0a0b:data=8'h00;
14'h0a0c:data=8'h00;
14'h0a0d:data=8'h00;
14'h0a0e:data=8'h00;
14'h0a0f:data=8'h00;
14'h0a10:data=8'h00;
14'h0a11:data=8'h00;
14'h0a12:data=8'h00;
14'h0a13:data=8'h00;
14'h0a14:data=8'h00;
14'h0a15:data=8'h00;
14'h0a16:data=8'h00;
14'h0a17:data=8'h00;
14'h0a18:data=8'h00;
14'h0a19:data=8'h07;
14'h0a1a:data=8'hFF;
14'h0a1b:data=8'hFF;
14'h0a1c:data=8'hFC;
14'h0a1d:data=8'h00;
14'h0a1e:data=8'h00;
14'h0a1f:data=8'h00;
14'h0a20:data=8'h00;
14'h0a21:data=8'h00;
14'h0a22:data=8'h1F;
14'h0a23:data=8'hFF;
14'h0a24:data=8'hFF;
14'h0a25:data=8'hFC;
14'h0a26:data=8'h00;
14'h0a27:data=8'h00;
14'h0a40:data=8'h01;
14'h0a41:data=8'hFF;
14'h0a42:data=8'hFF;
14'h0a43:data=8'hC0;
14'h0a44:data=8'h00;
14'h0a45:data=8'h00;
14'h0a46:data=8'h00;
14'h0a47:data=8'h00;
14'h0a48:data=8'h00;
14'h0a49:data=8'h00;
14'h0a4a:data=8'h00;
14'h0a4b:data=8'h00;
14'h0a4c:data=8'h00;
14'h0a4d:data=8'h00;
14'h0a4e:data=8'h00;
14'h0a4f:data=8'h00;
14'h0a50:data=8'h00;
14'h0a51:data=8'h00;
14'h0a52:data=8'h00;
14'h0a53:data=8'h00;
14'h0a54:data=8'h00;
14'h0a55:data=8'h00;
14'h0a56:data=8'h00;
14'h0a57:data=8'h00;
14'h0a58:data=8'h00;
14'h0a59:data=8'h07;
14'h0a5a:data=8'hFF;
14'h0a5b:data=8'hFF;
14'h0a5c:data=8'hFC;
14'h0a5d:data=8'h00;
14'h0a5e:data=8'h00;
14'h0a5f:data=8'h00;
14'h0a60:data=8'h00;
14'h0a61:data=8'h00;
14'h0a62:data=8'h1F;
14'h0a63:data=8'hFF;
14'h0a64:data=8'hFF;
14'h0a65:data=8'hFC;
14'h0a66:data=8'h00;
14'h0a67:data=8'h00;
14'h0a80:data=8'h01;
14'h0a81:data=8'hFF;
14'h0a82:data=8'hFF;
14'h0a83:data=8'hC0;
14'h0a84:data=8'h00;
14'h0a85:data=8'h00;
14'h0a86:data=8'h00;
14'h0a87:data=8'h00;
14'h0a88:data=8'h00;
14'h0a89:data=8'h00;
14'h0a8a:data=8'h00;
14'h0a8b:data=8'h00;
14'h0a8c:data=8'h00;
14'h0a8d:data=8'h00;
14'h0a8e:data=8'h00;
14'h0a8f:data=8'h00;
14'h0a90:data=8'h00;
14'h0a91:data=8'h00;
14'h0a92:data=8'h00;
14'h0a93:data=8'h00;
14'h0a94:data=8'h00;
14'h0a95:data=8'h00;
14'h0a96:data=8'h00;
14'h0a97:data=8'h00;
14'h0a98:data=8'h00;
14'h0a99:data=8'h07;
14'h0a9a:data=8'hFF;
14'h0a9b:data=8'hFF;
14'h0a9c:data=8'hFC;
14'h0a9d:data=8'h00;
14'h0a9e:data=8'h00;
14'h0a9f:data=8'h00;
14'h0aa0:data=8'h00;
14'h0aa1:data=8'h00;
14'h0aa2:data=8'h1F;
14'h0aa3:data=8'hFF;
14'h0aa4:data=8'hFF;
14'h0aa5:data=8'hFC;
14'h0aa6:data=8'h00;
14'h0aa7:data=8'h00;
14'h0ac0:data=8'h01;
14'h0ac1:data=8'hFF;
14'h0ac2:data=8'hFF;
14'h0ac3:data=8'hC0;
14'h0ac4:data=8'h00;
14'h0ac5:data=8'h00;
14'h0ac6:data=8'h00;
14'h0ac7:data=8'h00;
14'h0ac8:data=8'h00;
14'h0ac9:data=8'h00;
14'h0aca:data=8'h00;
14'h0acb:data=8'h00;
14'h0acc:data=8'h00;
14'h0acd:data=8'h00;
14'h0ace:data=8'h00;
14'h0acf:data=8'h00;
14'h0ad0:data=8'h00;
14'h0ad1:data=8'h00;
14'h0ad2:data=8'h00;
14'h0ad3:data=8'h00;
14'h0ad4:data=8'h00;
14'h0ad5:data=8'h00;
14'h0ad6:data=8'h00;
14'h0ad7:data=8'h00;
14'h0ad8:data=8'h00;
14'h0ad9:data=8'h07;
14'h0ada:data=8'hFF;
14'h0adb:data=8'hFF;
14'h0adc:data=8'hFC;
14'h0add:data=8'h00;
14'h0ade:data=8'h00;
14'h0adf:data=8'h00;
14'h0ae0:data=8'h00;
14'h0ae1:data=8'h00;
14'h0ae2:data=8'h1F;
14'h0ae3:data=8'hFF;
14'h0ae4:data=8'hFF;
14'h0ae5:data=8'hFC;
14'h0ae6:data=8'h00;
14'h0ae7:data=8'h00;
14'h0b00:data=8'h01;
14'h0b01:data=8'hFF;
14'h0b02:data=8'hFF;
14'h0b03:data=8'hC0;
14'h0b04:data=8'h00;
14'h0b05:data=8'h00;
14'h0b06:data=8'h00;
14'h0b07:data=8'h00;
14'h0b08:data=8'h00;
14'h0b09:data=8'h00;
14'h0b0a:data=8'h00;
14'h0b0b:data=8'h00;
14'h0b0c:data=8'h00;
14'h0b0d:data=8'h00;
14'h0b0e:data=8'h00;
14'h0b0f:data=8'h00;
14'h0b10:data=8'h00;
14'h0b11:data=8'h00;
14'h0b12:data=8'h00;
14'h0b13:data=8'h00;
14'h0b14:data=8'h00;
14'h0b15:data=8'h00;
14'h0b16:data=8'h00;
14'h0b17:data=8'h00;
14'h0b18:data=8'h00;
14'h0b19:data=8'h07;
14'h0b1a:data=8'hFF;
14'h0b1b:data=8'hFF;
14'h0b1c:data=8'hFC;
14'h0b1d:data=8'h00;
14'h0b1e:data=8'h00;
14'h0b1f:data=8'h00;
14'h0b20:data=8'h00;
14'h0b21:data=8'h00;
14'h0b22:data=8'h1F;
14'h0b23:data=8'hFF;
14'h0b24:data=8'hFF;
14'h0b25:data=8'hFC;
14'h0b26:data=8'h00;
14'h0b27:data=8'h00;
14'h0b40:data=8'h01;
14'h0b41:data=8'hFF;
14'h0b42:data=8'hFF;
14'h0b43:data=8'hC0;
14'h0b44:data=8'h00;
14'h0b45:data=8'h00;
14'h0b46:data=8'h00;
14'h0b47:data=8'h00;
14'h0b48:data=8'h00;
14'h0b49:data=8'h00;
14'h0b4a:data=8'h00;
14'h0b4b:data=8'h00;
14'h0b4c:data=8'h00;
14'h0b4d:data=8'h00;
14'h0b4e:data=8'h00;
14'h0b4f:data=8'h00;
14'h0b50:data=8'h00;
14'h0b51:data=8'h00;
14'h0b52:data=8'h00;
14'h0b53:data=8'h00;
14'h0b54:data=8'h00;
14'h0b55:data=8'h00;
14'h0b56:data=8'h00;
14'h0b57:data=8'h00;
14'h0b58:data=8'h00;
14'h0b59:data=8'h07;
14'h0b5a:data=8'hFF;
14'h0b5b:data=8'hFF;
14'h0b5c:data=8'hFC;
14'h0b5d:data=8'h00;
14'h0b5e:data=8'h00;
14'h0b5f:data=8'h00;
14'h0b60:data=8'h00;
14'h0b61:data=8'h00;
14'h0b62:data=8'h1F;
14'h0b63:data=8'hFF;
14'h0b64:data=8'hFF;
14'h0b65:data=8'hFC;
14'h0b66:data=8'h00;
14'h0b67:data=8'h00;
14'h0b80:data=8'h01;
14'h0b81:data=8'hFF;
14'h0b82:data=8'hFF;
14'h0b83:data=8'hC0;
14'h0b84:data=8'h00;
14'h0b85:data=8'h00;
14'h0b86:data=8'h00;
14'h0b87:data=8'h00;
14'h0b88:data=8'h00;
14'h0b89:data=8'h00;
14'h0b8a:data=8'h00;
14'h0b8b:data=8'h00;
14'h0b8c:data=8'h00;
14'h0b8d:data=8'h00;
14'h0b8e:data=8'h00;
14'h0b8f:data=8'h00;
14'h0b90:data=8'h00;
14'h0b91:data=8'h00;
14'h0b92:data=8'h00;
14'h0b93:data=8'h00;
14'h0b94:data=8'h00;
14'h0b95:data=8'h00;
14'h0b96:data=8'h00;
14'h0b97:data=8'h00;
14'h0b98:data=8'h00;
14'h0b99:data=8'h07;
14'h0b9a:data=8'hFF;
14'h0b9b:data=8'hFF;
14'h0b9c:data=8'hFC;
14'h0b9d:data=8'h00;
14'h0b9e:data=8'h00;
14'h0b9f:data=8'h00;
14'h0ba0:data=8'h00;
14'h0ba1:data=8'h00;
14'h0ba2:data=8'h1F;
14'h0ba3:data=8'hFF;
14'h0ba4:data=8'hFF;
14'h0ba5:data=8'hFC;
14'h0ba6:data=8'h00;
14'h0ba7:data=8'h00;
14'h0bc0:data=8'h01;
14'h0bc1:data=8'hFF;
14'h0bc2:data=8'hFF;
14'h0bc3:data=8'hC0;
14'h0bc4:data=8'h00;
14'h0bc5:data=8'h00;
14'h0bc6:data=8'h00;
14'h0bc7:data=8'h00;
14'h0bc8:data=8'h00;
14'h0bc9:data=8'h00;
14'h0bca:data=8'h00;
14'h0bcb:data=8'h00;
14'h0bcc:data=8'h00;
14'h0bcd:data=8'h00;
14'h0bce:data=8'h00;
14'h0bcf:data=8'h00;
14'h0bd0:data=8'h00;
14'h0bd1:data=8'h00;
14'h0bd2:data=8'h00;
14'h0bd3:data=8'h00;
14'h0bd4:data=8'h00;
14'h0bd5:data=8'h00;
14'h0bd6:data=8'h00;
14'h0bd7:data=8'h00;
14'h0bd8:data=8'h00;
14'h0bd9:data=8'h07;
14'h0bda:data=8'hFF;
14'h0bdb:data=8'hFF;
14'h0bdc:data=8'hFC;
14'h0bdd:data=8'h00;
14'h0bde:data=8'h00;
14'h0bdf:data=8'h00;
14'h0be0:data=8'h00;
14'h0be1:data=8'h00;
14'h0be2:data=8'h1F;
14'h0be3:data=8'hFF;
14'h0be4:data=8'hFF;
14'h0be5:data=8'hFC;
14'h0be6:data=8'h00;
14'h0be7:data=8'h00;
14'h0c00:data=8'h01;
14'h0c01:data=8'hFF;
14'h0c02:data=8'hFF;
14'h0c03:data=8'hC0;
14'h0c04:data=8'h00;
14'h0c05:data=8'h00;
14'h0c06:data=8'h00;
14'h0c07:data=8'h00;
14'h0c08:data=8'h00;
14'h0c09:data=8'h00;
14'h0c0a:data=8'h3F;
14'h0c0b:data=8'hE0;
14'h0c0c:data=8'h00;
14'h0c0d:data=8'h00;
14'h0c0e:data=8'h00;
14'h0c0f:data=8'h00;
14'h0c10:data=8'h00;
14'h0c11:data=8'h00;
14'h0c12:data=8'h00;
14'h0c13:data=8'h00;
14'h0c14:data=8'h00;
14'h0c15:data=8'h00;
14'h0c16:data=8'h00;
14'h0c17:data=8'h00;
14'h0c18:data=8'h00;
14'h0c19:data=8'h07;
14'h0c1a:data=8'hFF;
14'h0c1b:data=8'hFF;
14'h0c1c:data=8'hFC;
14'h0c1d:data=8'h00;
14'h0c1e:data=8'h00;
14'h0c1f:data=8'h00;
14'h0c20:data=8'h00;
14'h0c21:data=8'h00;
14'h0c22:data=8'h1F;
14'h0c23:data=8'hFF;
14'h0c24:data=8'hFF;
14'h0c25:data=8'hFC;
14'h0c26:data=8'h00;
14'h0c27:data=8'h00;
14'h0c40:data=8'h01;
14'h0c41:data=8'hFF;
14'h0c42:data=8'hFF;
14'h0c43:data=8'hC0;
14'h0c44:data=8'h00;
14'h0c45:data=8'h00;
14'h0c46:data=8'h00;
14'h0c47:data=8'h00;
14'h0c48:data=8'h00;
14'h0c49:data=8'h3F;
14'h0c4a:data=8'hFF;
14'h0c4b:data=8'hFE;
14'h0c4c:data=8'h00;
14'h0c4d:data=8'h00;
14'h0c4e:data=8'h00;
14'h0c4f:data=8'h00;
14'h0c50:data=8'h00;
14'h0c51:data=8'h00;
14'h0c52:data=8'h00;
14'h0c53:data=8'h00;
14'h0c54:data=8'h00;
14'h0c55:data=8'h00;
14'h0c56:data=8'h00;
14'h0c57:data=8'h00;
14'h0c58:data=8'h00;
14'h0c59:data=8'h07;
14'h0c5a:data=8'hFF;
14'h0c5b:data=8'hFF;
14'h0c5c:data=8'hFC;
14'h0c5d:data=8'h00;
14'h0c5e:data=8'h00;
14'h0c5f:data=8'h00;
14'h0c60:data=8'h00;
14'h0c61:data=8'h00;
14'h0c62:data=8'h1F;
14'h0c63:data=8'hFF;
14'h0c64:data=8'hFF;
14'h0c65:data=8'hFC;
14'h0c66:data=8'h00;
14'h0c67:data=8'h00;
14'h0c80:data=8'h01;
14'h0c81:data=8'hFF;
14'h0c82:data=8'hFF;
14'h0c83:data=8'hC0;
14'h0c84:data=8'h00;
14'h0c85:data=8'h00;
14'h0c86:data=8'h00;
14'h0c87:data=8'h00;
14'h0c88:data=8'h07;
14'h0c89:data=8'hFF;
14'h0c8a:data=8'hFF;
14'h0c8b:data=8'hFF;
14'h0c8c:data=8'hF0;
14'h0c8d:data=8'h00;
14'h0c8e:data=8'h00;
14'h0c8f:data=8'h00;
14'h0c90:data=8'h00;
14'h0c91:data=8'h00;
14'h0c92:data=8'h00;
14'h0c93:data=8'h00;
14'h0c94:data=8'h00;
14'h0c95:data=8'h00;
14'h0c96:data=8'h00;
14'h0c97:data=8'h00;
14'h0c98:data=8'h00;
14'h0c99:data=8'h07;
14'h0c9a:data=8'hFF;
14'h0c9b:data=8'hFF;
14'h0c9c:data=8'hFC;
14'h0c9d:data=8'h00;
14'h0c9e:data=8'h00;
14'h0c9f:data=8'h00;
14'h0ca0:data=8'h00;
14'h0ca1:data=8'h00;
14'h0ca2:data=8'h1F;
14'h0ca3:data=8'hFF;
14'h0ca4:data=8'hFF;
14'h0ca5:data=8'hFC;
14'h0ca6:data=8'h00;
14'h0ca7:data=8'h00;
14'h0cc0:data=8'h01;
14'h0cc1:data=8'hFF;
14'h0cc2:data=8'hFF;
14'h0cc3:data=8'hC0;
14'h0cc4:data=8'h00;
14'h0cc5:data=8'h00;
14'h0cc6:data=8'h00;
14'h0cc7:data=8'h00;
14'h0cc8:data=8'hFF;
14'h0cc9:data=8'hFF;
14'h0cca:data=8'hFF;
14'h0ccb:data=8'hFF;
14'h0ccc:data=8'hFE;
14'h0ccd:data=8'h00;
14'h0cce:data=8'h00;
14'h0ccf:data=8'h00;
14'h0cd0:data=8'h00;
14'h0cd1:data=8'h00;
14'h0cd2:data=8'h00;
14'h0cd3:data=8'h00;
14'h0cd4:data=8'h00;
14'h0cd5:data=8'h00;
14'h0cd6:data=8'h00;
14'h0cd7:data=8'h00;
14'h0cd8:data=8'h00;
14'h0cd9:data=8'h07;
14'h0cda:data=8'hFF;
14'h0cdb:data=8'hFF;
14'h0cdc:data=8'hFC;
14'h0cdd:data=8'h00;
14'h0cde:data=8'h00;
14'h0cdf:data=8'h00;
14'h0ce0:data=8'h00;
14'h0ce1:data=8'h00;
14'h0ce2:data=8'h1F;
14'h0ce3:data=8'hFF;
14'h0ce4:data=8'hFF;
14'h0ce5:data=8'hFC;
14'h0ce6:data=8'h00;
14'h0ce7:data=8'h00;
14'h0d00:data=8'h01;
14'h0d01:data=8'hFF;
14'h0d02:data=8'hFF;
14'h0d03:data=8'hC0;
14'h0d04:data=8'h00;
14'h0d05:data=8'h00;
14'h0d06:data=8'h00;
14'h0d07:data=8'h03;
14'h0d08:data=8'hFF;
14'h0d09:data=8'hFF;
14'h0d0a:data=8'hFF;
14'h0d0b:data=8'hFF;
14'h0d0c:data=8'hFF;
14'h0d0d:data=8'h80;
14'h0d0e:data=8'h00;
14'h0d0f:data=8'h00;
14'h0d10:data=8'h00;
14'h0d11:data=8'h00;
14'h0d12:data=8'h00;
14'h0d13:data=8'h00;
14'h0d14:data=8'h00;
14'h0d15:data=8'h00;
14'h0d16:data=8'h00;
14'h0d17:data=8'h00;
14'h0d18:data=8'h00;
14'h0d19:data=8'h07;
14'h0d1a:data=8'hFF;
14'h0d1b:data=8'hFF;
14'h0d1c:data=8'hFC;
14'h0d1d:data=8'h00;
14'h0d1e:data=8'h00;
14'h0d1f:data=8'h00;
14'h0d20:data=8'h00;
14'h0d21:data=8'h00;
14'h0d22:data=8'h1F;
14'h0d23:data=8'hFF;
14'h0d24:data=8'hFF;
14'h0d25:data=8'hFC;
14'h0d26:data=8'h00;
14'h0d27:data=8'h00;
14'h0d40:data=8'h01;
14'h0d41:data=8'hFF;
14'h0d42:data=8'hFF;
14'h0d43:data=8'hC0;
14'h0d44:data=8'h00;
14'h0d45:data=8'h00;
14'h0d46:data=8'h00;
14'h0d47:data=8'h1F;
14'h0d48:data=8'hFF;
14'h0d49:data=8'hFF;
14'h0d4a:data=8'hFF;
14'h0d4b:data=8'hFF;
14'h0d4c:data=8'hFF;
14'h0d4d:data=8'hF0;
14'h0d4e:data=8'h00;
14'h0d4f:data=8'h00;
14'h0d50:data=8'h00;
14'h0d51:data=8'h00;
14'h0d52:data=8'h00;
14'h0d53:data=8'h00;
14'h0d54:data=8'h00;
14'h0d55:data=8'h00;
14'h0d56:data=8'h00;
14'h0d57:data=8'h00;
14'h0d58:data=8'h00;
14'h0d59:data=8'h07;
14'h0d5a:data=8'hFF;
14'h0d5b:data=8'hFF;
14'h0d5c:data=8'hFC;
14'h0d5d:data=8'h00;
14'h0d5e:data=8'h00;
14'h0d5f:data=8'h00;
14'h0d60:data=8'h00;
14'h0d61:data=8'h00;
14'h0d62:data=8'h1F;
14'h0d63:data=8'hFF;
14'h0d64:data=8'hFF;
14'h0d65:data=8'hFC;
14'h0d66:data=8'h00;
14'h0d67:data=8'h00;
14'h0d80:data=8'h01;
14'h0d81:data=8'hFF;
14'h0d82:data=8'hFF;
14'h0d83:data=8'hC0;
14'h0d84:data=8'h00;
14'h0d85:data=8'h00;
14'h0d86:data=8'h00;
14'h0d87:data=8'hFF;
14'h0d88:data=8'hFF;
14'h0d89:data=8'hFF;
14'h0d8a:data=8'hFF;
14'h0d8b:data=8'hFF;
14'h0d8c:data=8'hFF;
14'h0d8d:data=8'hFC;
14'h0d8e:data=8'h00;
14'h0d8f:data=8'h00;
14'h0d90:data=8'h00;
14'h0d91:data=8'h00;
14'h0d92:data=8'h00;
14'h0d93:data=8'h00;
14'h0d94:data=8'h00;
14'h0d95:data=8'h00;
14'h0d96:data=8'h00;
14'h0d97:data=8'h00;
14'h0d98:data=8'h00;
14'h0d99:data=8'h07;
14'h0d9a:data=8'hFF;
14'h0d9b:data=8'hFF;
14'h0d9c:data=8'hFC;
14'h0d9d:data=8'h00;
14'h0d9e:data=8'h00;
14'h0d9f:data=8'h00;
14'h0da0:data=8'h00;
14'h0da1:data=8'h00;
14'h0da2:data=8'h1F;
14'h0da3:data=8'hFF;
14'h0da4:data=8'hFF;
14'h0da5:data=8'hFC;
14'h0da6:data=8'h00;
14'h0da7:data=8'h00;
14'h0dc0:data=8'h01;
14'h0dc1:data=8'hFF;
14'h0dc2:data=8'hFF;
14'h0dc3:data=8'hC0;
14'h0dc4:data=8'h00;
14'h0dc5:data=8'h00;
14'h0dc6:data=8'h03;
14'h0dc7:data=8'hFF;
14'h0dc8:data=8'hFF;
14'h0dc9:data=8'hFF;
14'h0dca:data=8'hFF;
14'h0dcb:data=8'hFF;
14'h0dcc:data=8'hFF;
14'h0dcd:data=8'hFF;
14'h0dce:data=8'h00;
14'h0dcf:data=8'h00;
14'h0dd0:data=8'h00;
14'h0dd1:data=8'h00;
14'h0dd2:data=8'h00;
14'h0dd3:data=8'h00;
14'h0dd4:data=8'h00;
14'h0dd5:data=8'h00;
14'h0dd6:data=8'h00;
14'h0dd7:data=8'h00;
14'h0dd8:data=8'h00;
14'h0dd9:data=8'h07;
14'h0dda:data=8'hFF;
14'h0ddb:data=8'hFF;
14'h0ddc:data=8'hFC;
14'h0ddd:data=8'h00;
14'h0dde:data=8'h00;
14'h0ddf:data=8'h00;
14'h0de0:data=8'h00;
14'h0de1:data=8'h00;
14'h0de2:data=8'h1F;
14'h0de3:data=8'hFF;
14'h0de4:data=8'hFF;
14'h0de5:data=8'hFC;
14'h0de6:data=8'h00;
14'h0de7:data=8'h00;
14'h0e00:data=8'h01;
14'h0e01:data=8'hFF;
14'h0e02:data=8'hFF;
14'h0e03:data=8'hC0;
14'h0e04:data=8'h00;
14'h0e05:data=8'h00;
14'h0e06:data=8'h0F;
14'h0e07:data=8'hFF;
14'h0e08:data=8'hFF;
14'h0e09:data=8'hFF;
14'h0e0a:data=8'hFF;
14'h0e0b:data=8'hFF;
14'h0e0c:data=8'hFF;
14'h0e0d:data=8'hFF;
14'h0e0e:data=8'hE0;
14'h0e0f:data=8'h00;
14'h0e10:data=8'h00;
14'h0e11:data=8'h00;
14'h0e12:data=8'h00;
14'h0e13:data=8'h00;
14'h0e14:data=8'h00;
14'h0e15:data=8'h00;
14'h0e16:data=8'h00;
14'h0e17:data=8'h00;
14'h0e18:data=8'h00;
14'h0e19:data=8'h07;
14'h0e1a:data=8'hFF;
14'h0e1b:data=8'hFF;
14'h0e1c:data=8'hFC;
14'h0e1d:data=8'h00;
14'h0e1e:data=8'h00;
14'h0e1f:data=8'h00;
14'h0e20:data=8'h00;
14'h0e21:data=8'h00;
14'h0e22:data=8'h1F;
14'h0e23:data=8'hFF;
14'h0e24:data=8'hFF;
14'h0e25:data=8'hFC;
14'h0e26:data=8'h00;
14'h0e27:data=8'h00;
14'h0e40:data=8'h01;
14'h0e41:data=8'hFF;
14'h0e42:data=8'hFF;
14'h0e43:data=8'hC0;
14'h0e44:data=8'h00;
14'h0e45:data=8'h00;
14'h0e46:data=8'h3F;
14'h0e47:data=8'hFF;
14'h0e48:data=8'hFF;
14'h0e49:data=8'hFF;
14'h0e4a:data=8'hFF;
14'h0e4b:data=8'hFF;
14'h0e4c:data=8'hFF;
14'h0e4d:data=8'hFF;
14'h0e4e:data=8'hF8;
14'h0e4f:data=8'h00;
14'h0e50:data=8'h00;
14'h0e51:data=8'h00;
14'h0e52:data=8'h00;
14'h0e53:data=8'h00;
14'h0e54:data=8'h00;
14'h0e55:data=8'h00;
14'h0e56:data=8'h00;
14'h0e57:data=8'h00;
14'h0e58:data=8'h00;
14'h0e59:data=8'h07;
14'h0e5a:data=8'hFF;
14'h0e5b:data=8'hFF;
14'h0e5c:data=8'hFC;
14'h0e5d:data=8'h00;
14'h0e5e:data=8'h00;
14'h0e5f:data=8'h00;
14'h0e60:data=8'h00;
14'h0e61:data=8'h00;
14'h0e62:data=8'h1F;
14'h0e63:data=8'hFF;
14'h0e64:data=8'hFF;
14'h0e65:data=8'hFC;
14'h0e66:data=8'h00;
14'h0e67:data=8'h00;
14'h0e80:data=8'h01;
14'h0e81:data=8'hFF;
14'h0e82:data=8'hFF;
14'h0e83:data=8'hC0;
14'h0e84:data=8'h00;
14'h0e85:data=8'h00;
14'h0e86:data=8'hFF;
14'h0e87:data=8'hFF;
14'h0e88:data=8'hFF;
14'h0e89:data=8'hFF;
14'h0e8a:data=8'hFF;
14'h0e8b:data=8'hFF;
14'h0e8c:data=8'hFF;
14'h0e8d:data=8'hFF;
14'h0e8e:data=8'hFF;
14'h0e8f:data=8'hC0;
14'h0e90:data=8'h00;
14'h0e91:data=8'h00;
14'h0e92:data=8'h00;
14'h0e93:data=8'h00;
14'h0e94:data=8'h00;
14'h0e95:data=8'h00;
14'h0e96:data=8'h00;
14'h0e97:data=8'h00;
14'h0e98:data=8'h00;
14'h0e99:data=8'h07;
14'h0e9a:data=8'hFF;
14'h0e9b:data=8'hFF;
14'h0e9c:data=8'hFC;
14'h0e9d:data=8'h00;
14'h0e9e:data=8'h00;
14'h0e9f:data=8'h00;
14'h0ea0:data=8'h00;
14'h0ea1:data=8'h00;
14'h0ea2:data=8'h1F;
14'h0ea3:data=8'hFF;
14'h0ea4:data=8'hFF;
14'h0ea5:data=8'hFC;
14'h0ea6:data=8'h00;
14'h0ea7:data=8'h00;
14'h0ec0:data=8'h01;
14'h0ec1:data=8'hFF;
14'h0ec2:data=8'hFF;
14'h0ec3:data=8'hC0;
14'h0ec4:data=8'h00;
14'h0ec5:data=8'h01;
14'h0ec6:data=8'hFF;
14'h0ec7:data=8'hFF;
14'h0ec8:data=8'hFF;
14'h0ec9:data=8'hFF;
14'h0eca:data=8'hFF;
14'h0ecb:data=8'hFF;
14'h0ecc:data=8'hFF;
14'h0ecd:data=8'hFF;
14'h0ece:data=8'hFF;
14'h0ecf:data=8'hFE;
14'h0ed0:data=8'h00;
14'h0ed1:data=8'h00;
14'h0ed2:data=8'h00;
14'h0ed3:data=8'h00;
14'h0ed4:data=8'h00;
14'h0ed5:data=8'h00;
14'h0ed6:data=8'h00;
14'h0ed7:data=8'h00;
14'h0ed8:data=8'h00;
14'h0ed9:data=8'h07;
14'h0eda:data=8'hFF;
14'h0edb:data=8'hFF;
14'h0edc:data=8'hFC;
14'h0edd:data=8'h00;
14'h0ede:data=8'h00;
14'h0edf:data=8'h00;
14'h0ee0:data=8'h00;
14'h0ee1:data=8'h00;
14'h0ee2:data=8'h1F;
14'h0ee3:data=8'hFF;
14'h0ee4:data=8'hFF;
14'h0ee5:data=8'hFC;
14'h0ee6:data=8'h00;
14'h0ee7:data=8'h00;
14'h0f00:data=8'h01;
14'h0f01:data=8'hFF;
14'h0f02:data=8'hFF;
14'h0f03:data=8'hC0;
14'h0f04:data=8'h00;
14'h0f05:data=8'h03;
14'h0f06:data=8'hFF;
14'h0f07:data=8'hFF;
14'h0f08:data=8'hFF;
14'h0f09:data=8'hFF;
14'h0f0a:data=8'hFF;
14'h0f0b:data=8'hFF;
14'h0f0c:data=8'hFF;
14'h0f0d:data=8'hFF;
14'h0f0e:data=8'hFF;
14'h0f0f:data=8'hFF;
14'h0f10:data=8'hF8;
14'h0f11:data=8'h00;
14'h0f12:data=8'h00;
14'h0f13:data=8'h00;
14'h0f14:data=8'h00;
14'h0f15:data=8'h00;
14'h0f16:data=8'h00;
14'h0f17:data=8'h00;
14'h0f18:data=8'h00;
14'h0f19:data=8'h07;
14'h0f1a:data=8'hFF;
14'h0f1b:data=8'hFF;
14'h0f1c:data=8'hFC;
14'h0f1d:data=8'h00;
14'h0f1e:data=8'h00;
14'h0f1f:data=8'h00;
14'h0f20:data=8'h00;
14'h0f21:data=8'h00;
14'h0f22:data=8'h1F;
14'h0f23:data=8'hFF;
14'h0f24:data=8'hFF;
14'h0f25:data=8'hFC;
14'h0f26:data=8'h00;
14'h0f27:data=8'h00;
14'h0f40:data=8'h01;
14'h0f41:data=8'hFF;
14'h0f42:data=8'hFF;
14'h0f43:data=8'hC0;
14'h0f44:data=8'h00;
14'h0f45:data=8'h07;
14'h0f46:data=8'hFF;
14'h0f47:data=8'hFF;
14'h0f48:data=8'hFF;
14'h0f49:data=8'hFF;
14'h0f4a:data=8'hFF;
14'h0f4b:data=8'hFF;
14'h0f4c:data=8'hFF;
14'h0f4d:data=8'hFF;
14'h0f4e:data=8'hFF;
14'h0f4f:data=8'hFF;
14'h0f50:data=8'hFF;
14'h0f51:data=8'hC0;
14'h0f52:data=8'h00;
14'h0f53:data=8'h00;
14'h0f54:data=8'h00;
14'h0f55:data=8'h00;
14'h0f56:data=8'h00;
14'h0f57:data=8'h00;
14'h0f58:data=8'h00;
14'h0f59:data=8'h07;
14'h0f5a:data=8'hFF;
14'h0f5b:data=8'hFF;
14'h0f5c:data=8'hFC;
14'h0f5d:data=8'h00;
14'h0f5e:data=8'h00;
14'h0f5f:data=8'h00;
14'h0f60:data=8'h00;
14'h0f61:data=8'h00;
14'h0f62:data=8'h1F;
14'h0f63:data=8'hFF;
14'h0f64:data=8'hFF;
14'h0f65:data=8'hFC;
14'h0f66:data=8'h00;
14'h0f67:data=8'h00;
14'h0f80:data=8'h01;
14'h0f81:data=8'hFF;
14'h0f82:data=8'hFF;
14'h0f83:data=8'hC0;
14'h0f84:data=8'h00;
14'h0f85:data=8'h0F;
14'h0f86:data=8'hFF;
14'h0f87:data=8'hFF;
14'h0f88:data=8'hFF;
14'h0f89:data=8'hFF;
14'h0f8a:data=8'hFF;
14'h0f8b:data=8'hFF;
14'h0f8c:data=8'hFF;
14'h0f8d:data=8'hFF;
14'h0f8e:data=8'hFF;
14'h0f8f:data=8'hFF;
14'h0f90:data=8'hFF;
14'h0f91:data=8'hFE;
14'h0f92:data=8'h00;
14'h0f93:data=8'h00;
14'h0f94:data=8'h00;
14'h0f95:data=8'h00;
14'h0f96:data=8'h00;
14'h0f97:data=8'h00;
14'h0f98:data=8'h00;
14'h0f99:data=8'h07;
14'h0f9a:data=8'hFF;
14'h0f9b:data=8'hFF;
14'h0f9c:data=8'hFC;
14'h0f9d:data=8'h00;
14'h0f9e:data=8'h00;
14'h0f9f:data=8'h00;
14'h0fa0:data=8'h00;
14'h0fa1:data=8'h00;
14'h0fa2:data=8'h1F;
14'h0fa3:data=8'hFF;
14'h0fa4:data=8'hFF;
14'h0fa5:data=8'hFC;
14'h0fa6:data=8'h00;
14'h0fa7:data=8'h00;
14'h0fc0:data=8'h01;
14'h0fc1:data=8'hFF;
14'h0fc2:data=8'hFF;
14'h0fc3:data=8'hC0;
14'h0fc4:data=8'h00;
14'h0fc5:data=8'h1F;
14'h0fc6:data=8'hFF;
14'h0fc7:data=8'hFF;
14'h0fc8:data=8'hFF;
14'h0fc9:data=8'hFF;
14'h0fca:data=8'hFF;
14'h0fcb:data=8'hFF;
14'h0fcc:data=8'hFF;
14'h0fcd:data=8'hFF;
14'h0fce:data=8'hFF;
14'h0fcf:data=8'hFF;
14'h0fd0:data=8'hFF;
14'h0fd1:data=8'hFF;
14'h0fd2:data=8'hF0;
14'h0fd3:data=8'h00;
14'h0fd4:data=8'h00;
14'h0fd5:data=8'h00;
14'h0fd6:data=8'h00;
14'h0fd7:data=8'h00;
14'h0fd8:data=8'h00;
14'h0fd9:data=8'h07;
14'h0fda:data=8'hFF;
14'h0fdb:data=8'hFF;
14'h0fdc:data=8'hFC;
14'h0fdd:data=8'h00;
14'h0fde:data=8'h00;
14'h0fdf:data=8'h00;
14'h0fe0:data=8'h00;
14'h0fe1:data=8'h00;
14'h0fe2:data=8'h1F;
14'h0fe3:data=8'hFF;
14'h0fe4:data=8'hFF;
14'h0fe5:data=8'hFC;
14'h0fe6:data=8'h00;
14'h0fe7:data=8'h00;
14'h1000:data=8'h01;
14'h1001:data=8'hFF;
14'h1002:data=8'hFF;
14'h1003:data=8'hC0;
14'h1004:data=8'h00;
14'h1005:data=8'h3F;
14'h1006:data=8'hFF;
14'h1007:data=8'hFF;
14'h1008:data=8'hFF;
14'h1009:data=8'hFF;
14'h100a:data=8'hFF;
14'h100b:data=8'hFF;
14'h100c:data=8'hFF;
14'h100d:data=8'hFF;
14'h100e:data=8'hFF;
14'h100f:data=8'hFF;
14'h1010:data=8'hFF;
14'h1011:data=8'hFF;
14'h1012:data=8'hFF;
14'h1013:data=8'hFF;
14'h1014:data=8'hFF;
14'h1015:data=8'hFF;
14'h1016:data=8'hE0;
14'h1017:data=8'h00;
14'h1018:data=8'h00;
14'h1019:data=8'h07;
14'h101a:data=8'hFF;
14'h101b:data=8'hFF;
14'h101c:data=8'hFC;
14'h101d:data=8'h00;
14'h101e:data=8'h00;
14'h101f:data=8'h00;
14'h1020:data=8'h00;
14'h1021:data=8'h00;
14'h1022:data=8'h1F;
14'h1023:data=8'hFF;
14'h1024:data=8'hFF;
14'h1025:data=8'hFC;
14'h1026:data=8'h00;
14'h1027:data=8'h00;
14'h1040:data=8'h01;
14'h1041:data=8'hFF;
14'h1042:data=8'hFF;
14'h1043:data=8'hC0;
14'h1044:data=8'h00;
14'h1045:data=8'h7F;
14'h1046:data=8'hFF;
14'h1047:data=8'hFF;
14'h1048:data=8'hFF;
14'h1049:data=8'hFF;
14'h104a:data=8'hFF;
14'h104b:data=8'hFF;
14'h104c:data=8'hFF;
14'h104d:data=8'hFF;
14'h104e:data=8'hFF;
14'h104f:data=8'hFF;
14'h1050:data=8'hFF;
14'h1051:data=8'hFF;
14'h1052:data=8'hFF;
14'h1053:data=8'hFF;
14'h1054:data=8'hFF;
14'h1055:data=8'hFF;
14'h1056:data=8'hE0;
14'h1057:data=8'h00;
14'h1058:data=8'h00;
14'h1059:data=8'h07;
14'h105a:data=8'hFF;
14'h105b:data=8'hFF;
14'h105c:data=8'hFC;
14'h105d:data=8'h00;
14'h105e:data=8'h00;
14'h105f:data=8'h00;
14'h1060:data=8'h00;
14'h1061:data=8'h00;
14'h1062:data=8'h1F;
14'h1063:data=8'hFF;
14'h1064:data=8'hC0;
14'h1065:data=8'h00;
14'h1066:data=8'h00;
14'h1067:data=8'h00;
14'h1080:data=8'h01;
14'h1081:data=8'hFF;
14'h1082:data=8'hFF;
14'h1083:data=8'hC0;
14'h1084:data=8'h00;
14'h1085:data=8'h7F;
14'h1086:data=8'hFF;
14'h1087:data=8'hFF;
14'h1088:data=8'hFF;
14'h1089:data=8'hFF;
14'h108a:data=8'hFF;
14'h108b:data=8'hFF;
14'h108c:data=8'hFF;
14'h108d:data=8'hFF;
14'h108e:data=8'hFF;
14'h108f:data=8'hFF;
14'h1090:data=8'hFF;
14'h1091:data=8'hFF;
14'h1092:data=8'hFF;
14'h1093:data=8'hFF;
14'h1094:data=8'hFF;
14'h1095:data=8'hFF;
14'h1096:data=8'hE0;
14'h1097:data=8'h00;
14'h1098:data=8'h00;
14'h1099:data=8'h07;
14'h109a:data=8'hFF;
14'h109b:data=8'hFF;
14'h109c:data=8'hFC;
14'h109d:data=8'h00;
14'h109e:data=8'h00;
14'h109f:data=8'h00;
14'h10a0:data=8'h00;
14'h10a1:data=8'h00;
14'h10a2:data=8'h00;
14'h10a3:data=8'h00;
14'h10a4:data=8'h00;
14'h10a5:data=8'h00;
14'h10a6:data=8'h00;
14'h10a7:data=8'h00;
14'h10c0:data=8'h01;
14'h10c1:data=8'hFF;
14'h10c2:data=8'hFF;
14'h10c3:data=8'hC0;
14'h10c4:data=8'h00;
14'h10c5:data=8'h7F;
14'h10c6:data=8'hFF;
14'h10c7:data=8'hFF;
14'h10c8:data=8'hFF;
14'h10c9:data=8'hFF;
14'h10ca:data=8'hFF;
14'h10cb:data=8'hFF;
14'h10cc:data=8'hFF;
14'h10cd:data=8'hFF;
14'h10ce:data=8'hFF;
14'h10cf:data=8'hFF;
14'h10d0:data=8'hFF;
14'h10d1:data=8'hFF;
14'h10d2:data=8'hFF;
14'h10d3:data=8'hFF;
14'h10d4:data=8'hFF;
14'h10d5:data=8'hFF;
14'h10d6:data=8'hE0;
14'h10d7:data=8'h00;
14'h10d8:data=8'h00;
14'h10d9:data=8'h07;
14'h10da:data=8'hFF;
14'h10db:data=8'hFF;
14'h10dc:data=8'hFC;
14'h10dd:data=8'h00;
14'h10de:data=8'h00;
14'h10df:data=8'h00;
14'h10e0:data=8'h00;
14'h10e1:data=8'h00;
14'h10e2:data=8'h00;
14'h10e3:data=8'h00;
14'h10e4:data=8'h00;
14'h10e5:data=8'h00;
14'h10e6:data=8'h00;
14'h10e7:data=8'h00;
14'h1100:data=8'h01;
14'h1101:data=8'hFF;
14'h1102:data=8'hFF;
14'h1103:data=8'hC0;
14'h1104:data=8'h00;
14'h1105:data=8'h7F;
14'h1106:data=8'hFF;
14'h1107:data=8'hFF;
14'h1108:data=8'hFF;
14'h1109:data=8'hFF;
14'h110a:data=8'hFF;
14'h110b:data=8'hFF;
14'h110c:data=8'hFF;
14'h110d:data=8'hFF;
14'h110e:data=8'hFF;
14'h110f:data=8'hFF;
14'h1110:data=8'hFF;
14'h1111:data=8'hFF;
14'h1112:data=8'hFF;
14'h1113:data=8'hFF;
14'h1114:data=8'hFF;
14'h1115:data=8'hFF;
14'h1116:data=8'hE0;
14'h1117:data=8'h00;
14'h1118:data=8'h00;
14'h1119:data=8'h00;
14'h111a:data=8'h00;
14'h111b:data=8'h00;
14'h111c:data=8'h00;
14'h111d:data=8'h00;
14'h111e:data=8'h00;
14'h111f:data=8'h00;
14'h1120:data=8'h00;
14'h1121:data=8'h00;
14'h1122:data=8'h00;
14'h1123:data=8'h00;
14'h1124:data=8'h00;
14'h1125:data=8'h00;
14'h1126:data=8'h00;
14'h1127:data=8'h00;
14'h1140:data=8'hFF;
14'h1141:data=8'hFF;
14'h1142:data=8'hFF;
14'h1143:data=8'hFF;
14'h1144:data=8'hFF;
14'h1145:data=8'hFF;
14'h1146:data=8'hFF;
14'h1147:data=8'hFF;
14'h1148:data=8'hFF;
14'h1149:data=8'hFF;
14'h114a:data=8'hFF;
14'h114b:data=8'hFF;
14'h114c:data=8'hFF;
14'h114d:data=8'hFF;
14'h114e:data=8'hFF;
14'h114f:data=8'hFF;
14'h1150:data=8'hFF;
14'h1151:data=8'hFF;
14'h1152:data=8'hFF;
14'h1153:data=8'hFF;
14'h1154:data=8'hFF;
14'h1155:data=8'hFF;
14'h1156:data=8'hFF;
14'h1157:data=8'hFF;
14'h1158:data=8'hFF;
14'h1159:data=8'hFF;
14'h115a:data=8'hFF;
14'h115b:data=8'hFF;
14'h115c:data=8'hFF;
14'h115d:data=8'hFF;
14'h115e:data=8'hFF;
14'h115f:data=8'hFF;
14'h1160:data=8'hFF;
14'h1161:data=8'hFF;
14'h1162:data=8'hFF;
14'h1163:data=8'hFF;
14'h1164:data=8'hFF;
14'h1165:data=8'hFF;
14'h1166:data=8'h00;
14'h1167:data=8'h00;
14'h1180:data=8'hFF;
14'h1181:data=8'hFF;
14'h1182:data=8'hFF;
14'h1183:data=8'hFF;
14'h1184:data=8'hFF;
14'h1185:data=8'hFF;
14'h1186:data=8'hFF;
14'h1187:data=8'hFF;
14'h1188:data=8'hFF;
14'h1189:data=8'hFF;
14'h118a:data=8'hFF;
14'h118b:data=8'hFF;
14'h118c:data=8'hFF;
14'h118d:data=8'hFF;
14'h118e:data=8'hFF;
14'h118f:data=8'hFF;
14'h1190:data=8'hFF;
14'h1191:data=8'hFF;
14'h1192:data=8'hFF;
14'h1193:data=8'hFF;
14'h1194:data=8'hFF;
14'h1195:data=8'hFF;
14'h1196:data=8'hFF;
14'h1197:data=8'hFF;
14'h1198:data=8'hFF;
14'h1199:data=8'hFF;
14'h119a:data=8'hFF;
14'h119b:data=8'hFF;
14'h119c:data=8'hFF;
14'h119d:data=8'hFF;
14'h119e:data=8'hFF;
14'h119f:data=8'hFF;
14'h11a0:data=8'hFF;
14'h11a1:data=8'hFF;
14'h11a2:data=8'hFF;
14'h11a3:data=8'hFF;
14'h11a4:data=8'hFF;
14'h11a5:data=8'hFF;
14'h11a6:data=8'h00;
14'h11a7:data=8'h00;
14'h11c0:data=8'hFF;
14'h11c1:data=8'hFF;
14'h11c2:data=8'hFF;
14'h11c3:data=8'hFF;
14'h11c4:data=8'hFF;
14'h11c5:data=8'hFF;
14'h11c6:data=8'hFF;
14'h11c7:data=8'hFF;
14'h11c8:data=8'hFF;
14'h11c9:data=8'hFF;
14'h11ca:data=8'hFF;
14'h11cb:data=8'hFF;
14'h11cc:data=8'hFF;
14'h11cd:data=8'hFF;
14'h11ce:data=8'hFF;
14'h11cf:data=8'hFF;
14'h11d0:data=8'hFF;
14'h11d1:data=8'hFF;
14'h11d2:data=8'hFF;
14'h11d3:data=8'hFF;
14'h11d4:data=8'hFF;
14'h11d5:data=8'hFF;
14'h11d6:data=8'hFF;
14'h11d7:data=8'hFF;
14'h11d8:data=8'hFF;
14'h11d9:data=8'hFF;
14'h11da:data=8'hFF;
14'h11db:data=8'hFF;
14'h11dc:data=8'hFF;
14'h11dd:data=8'hFF;
14'h11de:data=8'hFF;
14'h11df:data=8'hFF;
14'h11e0:data=8'hFF;
14'h11e1:data=8'hFF;
14'h11e2:data=8'hFF;
14'h11e3:data=8'hFF;
14'h11e4:data=8'hFF;
14'h11e5:data=8'hFF;
14'h11e6:data=8'h00;
14'h11e7:data=8'h00;
14'h1200:data=8'hFF;
14'h1201:data=8'hFF;
14'h1202:data=8'hFF;
14'h1203:data=8'hFF;
14'h1204:data=8'hFF;
14'h1205:data=8'hFF;
14'h1206:data=8'hFF;
14'h1207:data=8'hFF;
14'h1208:data=8'hFF;
14'h1209:data=8'hFF;
14'h120a:data=8'hFF;
14'h120b:data=8'hFF;
14'h120c:data=8'hFF;
14'h120d:data=8'hFF;
14'h120e:data=8'hFF;
14'h120f:data=8'hFF;
14'h1210:data=8'hFF;
14'h1211:data=8'hFF;
14'h1212:data=8'hFF;
14'h1213:data=8'hFF;
14'h1214:data=8'hFF;
14'h1215:data=8'hFF;
14'h1216:data=8'hFF;
14'h1217:data=8'hFF;
14'h1218:data=8'hFF;
14'h1219:data=8'hFF;
14'h121a:data=8'hFF;
14'h121b:data=8'hFF;
14'h121c:data=8'hFF;
14'h121d:data=8'hFF;
14'h121e:data=8'hFF;
14'h121f:data=8'hFF;
14'h1220:data=8'hFF;
14'h1221:data=8'hFF;
14'h1222:data=8'hFF;
14'h1223:data=8'hFF;
14'h1224:data=8'hFF;
14'h1225:data=8'hFF;
14'h1226:data=8'h00;
14'h1227:data=8'h00;
14'h1240:data=8'hFF;
14'h1241:data=8'hFF;
14'h1242:data=8'hFF;
14'h1243:data=8'hFF;
14'h1244:data=8'hFF;
14'h1245:data=8'hFF;
14'h1246:data=8'hFF;
14'h1247:data=8'hFF;
14'h1248:data=8'hFF;
14'h1249:data=8'hFF;
14'h124a:data=8'hFF;
14'h124b:data=8'hFF;
14'h124c:data=8'hFF;
14'h124d:data=8'hFF;
14'h124e:data=8'hFF;
14'h124f:data=8'hFF;
14'h1250:data=8'hFF;
14'h1251:data=8'hFF;
14'h1252:data=8'hFF;
14'h1253:data=8'hFF;
14'h1254:data=8'hFF;
14'h1255:data=8'hFF;
14'h1256:data=8'hFF;
14'h1257:data=8'hFF;
14'h1258:data=8'hFF;
14'h1259:data=8'hFF;
14'h125a:data=8'hFF;
14'h125b:data=8'hFF;
14'h125c:data=8'hFF;
14'h125d:data=8'hFF;
14'h125e:data=8'hFF;
14'h125f:data=8'hFF;
14'h1260:data=8'hFF;
14'h1261:data=8'hFF;
14'h1262:data=8'hFF;
14'h1263:data=8'hFF;
14'h1264:data=8'hFF;
14'h1265:data=8'hFF;
14'h1266:data=8'h00;
14'h1267:data=8'h00;
14'h1280:data=8'hFF;
14'h1281:data=8'hFF;
14'h1282:data=8'hFF;
14'h1283:data=8'hFF;
14'h1284:data=8'hFF;
14'h1285:data=8'hFF;
14'h1286:data=8'hFF;
14'h1287:data=8'hFF;
14'h1288:data=8'hFF;
14'h1289:data=8'hFF;
14'h128a:data=8'hFF;
14'h128b:data=8'hFF;
14'h128c:data=8'hFF;
14'h128d:data=8'hFF;
14'h128e:data=8'hFF;
14'h128f:data=8'hFF;
14'h1290:data=8'hFF;
14'h1291:data=8'hFF;
14'h1292:data=8'hFF;
14'h1293:data=8'hFF;
14'h1294:data=8'hFF;
14'h1295:data=8'hFF;
14'h1296:data=8'hFF;
14'h1297:data=8'hFF;
14'h1298:data=8'hFF;
14'h1299:data=8'hFF;
14'h129a:data=8'hFF;
14'h129b:data=8'hFF;
14'h129c:data=8'hFF;
14'h129d:data=8'hFF;
14'h129e:data=8'hFF;
14'h129f:data=8'hFF;
14'h12a0:data=8'hFF;
14'h12a1:data=8'hFF;
14'h12a2:data=8'hFF;
14'h12a3:data=8'hFF;
14'h12a4:data=8'hFF;
14'h12a5:data=8'hFF;
14'h12a6:data=8'h00;
14'h12a7:data=8'h00;
14'h12c0:data=8'hFF;
14'h12c1:data=8'hFF;
14'h12c2:data=8'hFF;
14'h12c3:data=8'hFF;
14'h12c4:data=8'hFF;
14'h12c5:data=8'hFF;
14'h12c6:data=8'hFF;
14'h12c7:data=8'hFF;
14'h12c8:data=8'hFF;
14'h12c9:data=8'hFF;
14'h12ca:data=8'hFF;
14'h12cb:data=8'hFF;
14'h12cc:data=8'hFF;
14'h12cd:data=8'hFF;
14'h12ce:data=8'hFF;
14'h12cf:data=8'hFF;
14'h12d0:data=8'hFF;
14'h12d1:data=8'hFF;
14'h12d2:data=8'hFF;
14'h12d3:data=8'hFF;
14'h12d4:data=8'hFF;
14'h12d5:data=8'hFF;
14'h12d6:data=8'hFF;
14'h12d7:data=8'hFF;
14'h12d8:data=8'hFF;
14'h12d9:data=8'hFF;
14'h12da:data=8'hFF;
14'h12db:data=8'hFF;
14'h12dc:data=8'hFF;
14'h12dd:data=8'hFF;
14'h12de:data=8'hFF;
14'h12df:data=8'hFF;
14'h12e0:data=8'hFF;
14'h12e1:data=8'hFF;
14'h12e2:data=8'hFF;
14'h12e3:data=8'hFF;
14'h12e4:data=8'hFF;
14'h12e5:data=8'hFF;
14'h12e6:data=8'h00;
14'h12e7:data=8'h00;
14'h1300:data=8'hFF;
14'h1301:data=8'hFF;
14'h1302:data=8'hFF;
14'h1303:data=8'hFF;
14'h1304:data=8'hFF;
14'h1305:data=8'hFF;
14'h1306:data=8'hFF;
14'h1307:data=8'hFF;
14'h1308:data=8'hFF;
14'h1309:data=8'hFF;
14'h130a:data=8'hFF;
14'h130b:data=8'hFF;
14'h130c:data=8'hFF;
14'h130d:data=8'hFF;
14'h130e:data=8'hFF;
14'h130f:data=8'hFF;
14'h1310:data=8'hFF;
14'h1311:data=8'hFF;
14'h1312:data=8'hFF;
14'h1313:data=8'hFF;
14'h1314:data=8'hFF;
14'h1315:data=8'hFF;
14'h1316:data=8'hFF;
14'h1317:data=8'hFF;
14'h1318:data=8'hFF;
14'h1319:data=8'hFF;
14'h131a:data=8'hFF;
14'h131b:data=8'hFF;
14'h131c:data=8'hFF;
14'h131d:data=8'hFF;
14'h131e:data=8'hFF;
14'h131f:data=8'hFF;
14'h1320:data=8'hFF;
14'h1321:data=8'hFF;
14'h1322:data=8'hFF;
14'h1323:data=8'hFF;
14'h1324:data=8'hFF;
14'h1325:data=8'hFF;
14'h1326:data=8'h00;
14'h1327:data=8'h00;
14'h1340:data=8'hFF;
14'h1341:data=8'hFF;
14'h1342:data=8'hFF;
14'h1343:data=8'hFF;
14'h1344:data=8'hFF;
14'h1345:data=8'hFF;
14'h1346:data=8'hFF;
14'h1347:data=8'hFF;
14'h1348:data=8'hFF;
14'h1349:data=8'hFF;
14'h134a:data=8'hFF;
14'h134b:data=8'hFF;
14'h134c:data=8'hFF;
14'h134d:data=8'hFF;
14'h134e:data=8'hFF;
14'h134f:data=8'hFF;
14'h1350:data=8'hFF;
14'h1351:data=8'hFF;
14'h1352:data=8'hFF;
14'h1353:data=8'hFF;
14'h1354:data=8'hFF;
14'h1355:data=8'hFF;
14'h1356:data=8'hFF;
14'h1357:data=8'hFF;
14'h1358:data=8'hFF;
14'h1359:data=8'hFF;
14'h135a:data=8'hFF;
14'h135b:data=8'hFF;
14'h135c:data=8'hFF;
14'h135d:data=8'hFF;
14'h135e:data=8'hFF;
14'h135f:data=8'hFF;
14'h1360:data=8'hFF;
14'h1361:data=8'hFF;
14'h1362:data=8'hFF;
14'h1363:data=8'hFF;
14'h1364:data=8'hFF;
14'h1365:data=8'hFF;
14'h1366:data=8'h00;
14'h1367:data=8'h00;
14'h1380:data=8'hFF;
14'h1381:data=8'hFF;
14'h1382:data=8'hFF;
14'h1383:data=8'hFF;
14'h1384:data=8'hFF;
14'h1385:data=8'hFF;
14'h1386:data=8'hFF;
14'h1387:data=8'hFF;
14'h1388:data=8'hFF;
14'h1389:data=8'hFF;
14'h138a:data=8'hFF;
14'h138b:data=8'hFF;
14'h138c:data=8'hFF;
14'h138d:data=8'hFF;
14'h138e:data=8'hFF;
14'h138f:data=8'hFF;
14'h1390:data=8'hFF;
14'h1391:data=8'hFF;
14'h1392:data=8'hFF;
14'h1393:data=8'hFF;
14'h1394:data=8'hFF;
14'h1395:data=8'hFF;
14'h1396:data=8'hFF;
14'h1397:data=8'hFF;
14'h1398:data=8'hFF;
14'h1399:data=8'hFF;
14'h139a:data=8'hFF;
14'h139b:data=8'hFF;
14'h139c:data=8'hFF;
14'h139d:data=8'hFF;
14'h139e:data=8'hFF;
14'h139f:data=8'hFF;
14'h13a0:data=8'hFF;
14'h13a1:data=8'hFF;
14'h13a2:data=8'hFF;
14'h13a3:data=8'hFF;
14'h13a4:data=8'hFF;
14'h13a5:data=8'hFF;
14'h13a6:data=8'h00;
14'h13a7:data=8'h00;
14'h13c0:data=8'hFF;
14'h13c1:data=8'hFF;
14'h13c2:data=8'hFF;
14'h13c3:data=8'hFF;
14'h13c4:data=8'hFF;
14'h13c5:data=8'hFF;
14'h13c6:data=8'hFF;
14'h13c7:data=8'hFF;
14'h13c8:data=8'hFF;
14'h13c9:data=8'hFF;
14'h13ca:data=8'hFF;
14'h13cb:data=8'hFF;
14'h13cc:data=8'hFF;
14'h13cd:data=8'hFF;
14'h13ce:data=8'hFF;
14'h13cf:data=8'hFF;
14'h13d0:data=8'hFF;
14'h13d1:data=8'hFF;
14'h13d2:data=8'hFF;
14'h13d3:data=8'hFF;
14'h13d4:data=8'hFF;
14'h13d5:data=8'hFF;
14'h13d6:data=8'hFF;
14'h13d7:data=8'hFF;
14'h13d8:data=8'hFF;
14'h13d9:data=8'hFF;
14'h13da:data=8'hFF;
14'h13db:data=8'hFF;
14'h13dc:data=8'hFF;
14'h13dd:data=8'hFF;
14'h13de:data=8'hFF;
14'h13df:data=8'hFF;
14'h13e0:data=8'hFF;
14'h13e1:data=8'hFF;
14'h13e2:data=8'hFF;
14'h13e3:data=8'hFF;
14'h13e4:data=8'hFF;
14'h13e5:data=8'hFF;
14'h13e6:data=8'h00;
14'h13e7:data=8'h00;
14'h1400:data=8'hFF;
14'h1401:data=8'hFF;
14'h1402:data=8'hFF;
14'h1403:data=8'hFF;
14'h1404:data=8'hFF;
14'h1405:data=8'hFF;
14'h1406:data=8'hFF;
14'h1407:data=8'hFF;
14'h1408:data=8'hFF;
14'h1409:data=8'hFF;
14'h140a:data=8'hFF;
14'h140b:data=8'hFF;
14'h140c:data=8'hFF;
14'h140d:data=8'hFF;
14'h140e:data=8'hFF;
14'h140f:data=8'hFF;
14'h1410:data=8'hFF;
14'h1411:data=8'hFF;
14'h1412:data=8'hFF;
14'h1413:data=8'hFF;
14'h1414:data=8'hFF;
14'h1415:data=8'hFF;
14'h1416:data=8'hFF;
14'h1417:data=8'hFF;
14'h1418:data=8'hFF;
14'h1419:data=8'hFF;
14'h141a:data=8'hFF;
14'h141b:data=8'hFF;
14'h141c:data=8'hFF;
14'h141d:data=8'hFF;
14'h141e:data=8'hFF;
14'h141f:data=8'hFF;
14'h1420:data=8'hFF;
14'h1421:data=8'hFF;
14'h1422:data=8'hFF;
14'h1423:data=8'hFF;
14'h1424:data=8'hFF;
14'h1425:data=8'hFF;
14'h1426:data=8'h00;
14'h1427:data=8'h00;
14'h1440:data=8'hFF;
14'h1441:data=8'hFF;
14'h1442:data=8'hFF;
14'h1443:data=8'hFF;
14'h1444:data=8'hFF;
14'h1445:data=8'hFF;
14'h1446:data=8'hFF;
14'h1447:data=8'hFF;
14'h1448:data=8'hFF;
14'h1449:data=8'hFF;
14'h144a:data=8'hFF;
14'h144b:data=8'hFF;
14'h144c:data=8'hFF;
14'h144d:data=8'hFF;
14'h144e:data=8'hFF;
14'h144f:data=8'hFF;
14'h1450:data=8'hFF;
14'h1451:data=8'hFF;
14'h1452:data=8'hFF;
14'h1453:data=8'hFF;
14'h1454:data=8'hFF;
14'h1455:data=8'hFF;
14'h1456:data=8'hFF;
14'h1457:data=8'hFF;
14'h1458:data=8'hFF;
14'h1459:data=8'hFF;
14'h145a:data=8'hFF;
14'h145b:data=8'hFF;
14'h145c:data=8'hFF;
14'h145d:data=8'hFF;
14'h145e:data=8'hFF;
14'h145f:data=8'hFF;
14'h1460:data=8'hFF;
14'h1461:data=8'hFF;
14'h1462:data=8'hFF;
14'h1463:data=8'hFF;
14'h1464:data=8'hFF;
14'h1465:data=8'hFF;
14'h1466:data=8'h00;
14'h1467:data=8'h00;
14'h1480:data=8'hFF;
14'h1481:data=8'hFF;
14'h1482:data=8'hFF;
14'h1483:data=8'hFF;
14'h1484:data=8'hFF;
14'h1485:data=8'hFF;
14'h1486:data=8'hFF;
14'h1487:data=8'hFF;
14'h1488:data=8'hFF;
14'h1489:data=8'hFF;
14'h148a:data=8'hFF;
14'h148b:data=8'hFF;
14'h148c:data=8'hFF;
14'h148d:data=8'hFF;
14'h148e:data=8'hFF;
14'h148f:data=8'hFF;
14'h1490:data=8'hFF;
14'h1491:data=8'hFF;
14'h1492:data=8'hFF;
14'h1493:data=8'hFF;
14'h1494:data=8'hFF;
14'h1495:data=8'hFF;
14'h1496:data=8'hFF;
14'h1497:data=8'hFF;
14'h1498:data=8'hFF;
14'h1499:data=8'hFF;
14'h149a:data=8'hFF;
14'h149b:data=8'hFF;
14'h149c:data=8'hFF;
14'h149d:data=8'hFF;
14'h149e:data=8'hFF;
14'h149f:data=8'hFF;
14'h14a0:data=8'hFF;
14'h14a1:data=8'hFF;
14'h14a2:data=8'hFF;
14'h14a3:data=8'hFF;
14'h14a4:data=8'hFF;
14'h14a5:data=8'hFF;
14'h14a6:data=8'h00;
14'h14a7:data=8'h00;
14'h14c0:data=8'hFF;
14'h14c1:data=8'hFF;
14'h14c2:data=8'hFF;
14'h14c3:data=8'hFF;
14'h14c4:data=8'hFF;
14'h14c5:data=8'hFF;
14'h14c6:data=8'hFF;
14'h14c7:data=8'hFF;
14'h14c8:data=8'hFF;
14'h14c9:data=8'hFF;
14'h14ca:data=8'hFF;
14'h14cb:data=8'hFF;
14'h14cc:data=8'hFF;
14'h14cd:data=8'hFF;
14'h14ce:data=8'hFF;
14'h14cf:data=8'hFF;
14'h14d0:data=8'hFF;
14'h14d1:data=8'hFF;
14'h14d2:data=8'hFF;
14'h14d3:data=8'hFF;
14'h14d4:data=8'hFF;
14'h14d5:data=8'hFF;
14'h14d6:data=8'hFF;
14'h14d7:data=8'hFF;
14'h14d8:data=8'hFF;
14'h14d9:data=8'hFF;
14'h14da:data=8'hFF;
14'h14db:data=8'hFF;
14'h14dc:data=8'hFF;
14'h14dd:data=8'hFF;
14'h14de:data=8'hFF;
14'h14df:data=8'hFF;
14'h14e0:data=8'hFF;
14'h14e1:data=8'hFF;
14'h14e2:data=8'hFF;
14'h14e3:data=8'hFF;
14'h14e4:data=8'hFF;
14'h14e5:data=8'hFF;
14'h14e6:data=8'h00;
14'h14e7:data=8'h00;
14'h1500:data=8'hFF;
14'h1501:data=8'hFF;
14'h1502:data=8'hFF;
14'h1503:data=8'hFF;
14'h1504:data=8'hFF;
14'h1505:data=8'hFF;
14'h1506:data=8'hFF;
14'h1507:data=8'hFF;
14'h1508:data=8'hFF;
14'h1509:data=8'hFF;
14'h150a:data=8'hFF;
14'h150b:data=8'hFF;
14'h150c:data=8'hFF;
14'h150d:data=8'hFF;
14'h150e:data=8'hFF;
14'h150f:data=8'hFF;
14'h1510:data=8'hFF;
14'h1511:data=8'hFF;
14'h1512:data=8'hFF;
14'h1513:data=8'hFF;
14'h1514:data=8'hFF;
14'h1515:data=8'hFF;
14'h1516:data=8'hFF;
14'h1517:data=8'hFF;
14'h1518:data=8'hFF;
14'h1519:data=8'hFF;
14'h151a:data=8'hFF;
14'h151b:data=8'hFF;
14'h151c:data=8'hFF;
14'h151d:data=8'hFF;
14'h151e:data=8'hFF;
14'h151f:data=8'hFF;
14'h1520:data=8'hFF;
14'h1521:data=8'hFF;
14'h1522:data=8'hFF;
14'h1523:data=8'hFF;
14'h1524:data=8'hFF;
14'h1525:data=8'hFF;
14'h1526:data=8'h00;
14'h1527:data=8'h00;
14'h1540:data=8'h00;
14'h1541:data=8'h00;
14'h1542:data=8'h00;
14'h1543:data=8'h00;
14'h1544:data=8'h00;
14'h1545:data=8'h00;
14'h1546:data=8'h00;
14'h1547:data=8'h00;
14'h1548:data=8'h00;
14'h1549:data=8'h00;
14'h154a:data=8'h00;
14'h154b:data=8'h00;
14'h154c:data=8'h00;
14'h154d:data=8'h00;
14'h154e:data=8'h00;
14'h154f:data=8'h00;
14'h1550:data=8'h00;
14'h1551:data=8'h00;
14'h1552:data=8'h00;
14'h1553:data=8'h00;
14'h1554:data=8'h00;
14'h1555:data=8'h00;
14'h1556:data=8'h00;
14'h1557:data=8'h00;
14'h1558:data=8'h00;
14'h1559:data=8'h00;
14'h155a:data=8'h00;
14'h155b:data=8'h00;
14'h155c:data=8'h00;
14'h155d:data=8'h00;
14'h155e:data=8'h00;
14'h155f:data=8'h00;
14'h1560:data=8'h00;
14'h1561:data=8'h00;
14'h1562:data=8'h00;
14'h1563:data=8'h00;
14'h1564:data=8'h00;
14'h1565:data=8'h00;
14'h1566:data=8'h00;
14'h1567:data=8'h00;
14'h1580:data=8'h00;
14'h1581:data=8'h00;
14'h1582:data=8'h00;
14'h1583:data=8'h00;
14'h1584:data=8'h00;
14'h1585:data=8'h00;
14'h1586:data=8'h00;
14'h1587:data=8'h00;
14'h1588:data=8'h00;
14'h1589:data=8'h00;
14'h158a:data=8'h00;
14'h158b:data=8'h00;
14'h158c:data=8'h00;
14'h158d:data=8'h00;
14'h158e:data=8'h00;
14'h158f:data=8'h00;
14'h1590:data=8'h00;
14'h1591:data=8'h00;
14'h1592:data=8'h00;
14'h1593:data=8'h00;
14'h1594:data=8'h00;
14'h1595:data=8'h00;
14'h1596:data=8'h00;
14'h1597:data=8'h00;
14'h1598:data=8'h00;
14'h1599:data=8'h00;
14'h159a:data=8'h00;
14'h159b:data=8'h00;
14'h159c:data=8'h00;
14'h159d:data=8'h00;
14'h159e:data=8'h00;
14'h159f:data=8'h00;
14'h15a0:data=8'h00;
14'h15a1:data=8'h00;
14'h15a2:data=8'h00;
14'h15a3:data=8'h00;
14'h15a4:data=8'h00;
14'h15a5:data=8'h00;
14'h15a6:data=8'h00;
14'h15a7:data=8'h00;
14'h15c0:data=8'h00;
14'h15c1:data=8'h00;
14'h15c2:data=8'h00;
14'h15c3:data=8'h00;
14'h15c4:data=8'h00;
14'h15c5:data=8'h00;
14'h15c6:data=8'h00;
14'h15c7:data=8'h00;
14'h15c8:data=8'h00;
14'h15c9:data=8'h00;
14'h15ca:data=8'h00;
14'h15cb:data=8'h00;
14'h15cc:data=8'h00;
14'h15cd:data=8'h00;
14'h15ce:data=8'h00;
14'h15cf:data=8'h00;
14'h15d0:data=8'h00;
14'h15d1:data=8'h07;
14'h15d2:data=8'hFF;
14'h15d3:data=8'hFE;
14'h15d4:data=8'h00;
14'h15d5:data=8'h00;
14'h15d6:data=8'h00;
14'h15d7:data=8'h00;
14'h15d8:data=8'h00;
14'h15d9:data=8'h00;
14'h15da:data=8'h00;
14'h15db:data=8'h00;
14'h15dc:data=8'h00;
14'h15dd:data=8'h00;
14'h15de:data=8'h00;
14'h15df:data=8'h00;
14'h15e0:data=8'h00;
14'h15e1:data=8'h00;
14'h15e2:data=8'h00;
14'h15e3:data=8'h00;
14'h15e4:data=8'h00;
14'h15e5:data=8'h00;
14'h15e6:data=8'h00;
14'h15e7:data=8'h00;
14'h1600:data=8'h00;
14'h1601:data=8'h00;
14'h1602:data=8'h00;
14'h1603:data=8'h00;
14'h1604:data=8'h00;
14'h1605:data=8'h00;
14'h1606:data=8'h00;
14'h1607:data=8'h00;
14'h1608:data=8'h00;
14'h1609:data=8'h00;
14'h160a:data=8'h00;
14'h160b:data=8'h00;
14'h160c:data=8'h00;
14'h160d:data=8'h00;
14'h160e:data=8'h00;
14'h160f:data=8'h00;
14'h1610:data=8'h00;
14'h1611:data=8'h07;
14'h1612:data=8'hFF;
14'h1613:data=8'hFE;
14'h1614:data=8'h00;
14'h1615:data=8'h00;
14'h1616:data=8'h00;
14'h1617:data=8'h00;
14'h1618:data=8'h00;
14'h1619:data=8'h00;
14'h161a:data=8'h00;
14'h161b:data=8'h00;
14'h161c:data=8'h00;
14'h161d:data=8'h00;
14'h161e:data=8'h00;
14'h161f:data=8'h00;
14'h1620:data=8'h00;
14'h1621:data=8'h00;
14'h1622:data=8'h00;
14'h1623:data=8'h00;
14'h1624:data=8'h00;
14'h1625:data=8'h00;
14'h1626:data=8'h00;
14'h1627:data=8'h00;
14'h1640:data=8'h00;
14'h1641:data=8'h00;
14'h1642:data=8'h00;
14'h1643:data=8'h00;
14'h1644:data=8'h00;
14'h1645:data=8'h00;
14'h1646:data=8'h00;
14'h1647:data=8'h00;
14'h1648:data=8'h00;
14'h1649:data=8'h00;
14'h164a:data=8'h07;
14'h164b:data=8'hFF;
14'h164c:data=8'hF8;
14'h164d:data=8'h00;
14'h164e:data=8'h00;
14'h164f:data=8'h00;
14'h1650:data=8'h00;
14'h1651:data=8'h07;
14'h1652:data=8'hFF;
14'h1653:data=8'hFE;
14'h1654:data=8'h00;
14'h1655:data=8'h00;
14'h1656:data=8'h00;
14'h1657:data=8'h00;
14'h1658:data=8'h00;
14'h1659:data=8'h00;
14'h165a:data=8'h00;
14'h165b:data=8'h00;
14'h165c:data=8'h00;
14'h165d:data=8'h00;
14'h165e:data=8'h00;
14'h165f:data=8'h00;
14'h1660:data=8'h00;
14'h1661:data=8'h00;
14'h1662:data=8'h00;
14'h1663:data=8'h00;
14'h1664:data=8'h00;
14'h1665:data=8'h00;
14'h1666:data=8'h00;
14'h1667:data=8'h00;
14'h1680:data=8'h00;
14'h1681:data=8'h00;
14'h1682:data=8'h00;
14'h1683:data=8'h00;
14'h1684:data=8'h00;
14'h1685:data=8'h00;
14'h1686:data=8'h00;
14'h1687:data=8'h00;
14'h1688:data=8'h00;
14'h1689:data=8'h00;
14'h168a:data=8'h07;
14'h168b:data=8'hFF;
14'h168c:data=8'hF8;
14'h168d:data=8'h00;
14'h168e:data=8'h00;
14'h168f:data=8'h00;
14'h1690:data=8'h00;
14'h1691:data=8'h07;
14'h1692:data=8'hFF;
14'h1693:data=8'hFE;
14'h1694:data=8'h00;
14'h1695:data=8'h00;
14'h1696:data=8'h00;
14'h1697:data=8'h00;
14'h1698:data=8'h00;
14'h1699:data=8'h00;
14'h169a:data=8'h00;
14'h169b:data=8'h00;
14'h169c:data=8'h00;
14'h169d:data=8'h00;
14'h169e:data=8'h00;
14'h169f:data=8'h00;
14'h16a0:data=8'h00;
14'h16a1:data=8'h00;
14'h16a2:data=8'h00;
14'h16a3:data=8'h00;
14'h16a4:data=8'h00;
14'h16a5:data=8'h00;
14'h16a6:data=8'h00;
14'h16a7:data=8'h00;
14'h16c0:data=8'h00;
14'h16c1:data=8'h00;
14'h16c2:data=8'h00;
14'h16c3:data=8'h00;
14'h16c4:data=8'h00;
14'h16c5:data=8'h00;
14'h16c6:data=8'h00;
14'h16c7:data=8'h00;
14'h16c8:data=8'h00;
14'h16c9:data=8'h00;
14'h16ca:data=8'h07;
14'h16cb:data=8'hFF;
14'h16cc:data=8'hF8;
14'h16cd:data=8'h00;
14'h16ce:data=8'h00;
14'h16cf:data=8'h00;
14'h16d0:data=8'h00;
14'h16d1:data=8'h07;
14'h16d2:data=8'hFF;
14'h16d3:data=8'hFE;
14'h16d4:data=8'h00;
14'h16d5:data=8'h00;
14'h16d6:data=8'h00;
14'h16d7:data=8'h00;
14'h16d8:data=8'h00;
14'h16d9:data=8'h00;
14'h16da:data=8'h00;
14'h16db:data=8'h00;
14'h16dc:data=8'h00;
14'h16dd:data=8'h00;
14'h16de:data=8'h00;
14'h16df:data=8'h00;
14'h16e0:data=8'h00;
14'h16e1:data=8'h00;
14'h16e2:data=8'h00;
14'h16e3:data=8'h00;
14'h16e4:data=8'h00;
14'h16e5:data=8'h00;
14'h16e6:data=8'h00;
14'h16e7:data=8'h00;
14'h1700:data=8'h00;
14'h1701:data=8'h00;
14'h1702:data=8'h00;
14'h1703:data=8'h00;
14'h1704:data=8'h00;
14'h1705:data=8'h00;
14'h1706:data=8'h00;
14'h1707:data=8'h00;
14'h1708:data=8'h00;
14'h1709:data=8'h00;
14'h170a:data=8'h07;
14'h170b:data=8'hFF;
14'h170c:data=8'hF8;
14'h170d:data=8'h00;
14'h170e:data=8'h00;
14'h170f:data=8'h00;
14'h1710:data=8'h00;
14'h1711:data=8'h07;
14'h1712:data=8'hFF;
14'h1713:data=8'hFE;
14'h1714:data=8'h00;
14'h1715:data=8'h00;
14'h1716:data=8'h00;
14'h1717:data=8'h00;
14'h1718:data=8'h00;
14'h1719:data=8'h00;
14'h171a:data=8'h00;
14'h171b:data=8'h00;
14'h171c:data=8'h00;
14'h171d:data=8'h00;
14'h171e:data=8'h00;
14'h171f:data=8'h00;
14'h1720:data=8'h00;
14'h1721:data=8'h00;
14'h1722:data=8'h00;
14'h1723:data=8'h00;
14'h1724:data=8'h00;
14'h1725:data=8'h00;
14'h1726:data=8'h00;
14'h1727:data=8'h00;
14'h1740:data=8'h00;
14'h1741:data=8'h00;
14'h1742:data=8'h00;
14'h1743:data=8'h00;
14'h1744:data=8'h00;
14'h1745:data=8'h00;
14'h1746:data=8'h00;
14'h1747:data=8'h00;
14'h1748:data=8'h00;
14'h1749:data=8'h00;
14'h174a:data=8'h07;
14'h174b:data=8'hFF;
14'h174c:data=8'hF8;
14'h174d:data=8'h00;
14'h174e:data=8'h00;
14'h174f:data=8'h00;
14'h1750:data=8'h00;
14'h1751:data=8'h07;
14'h1752:data=8'hFF;
14'h1753:data=8'hFE;
14'h1754:data=8'h00;
14'h1755:data=8'h00;
14'h1756:data=8'h00;
14'h1757:data=8'h00;
14'h1758:data=8'h00;
14'h1759:data=8'h00;
14'h175a:data=8'h00;
14'h175b:data=8'h00;
14'h175c:data=8'h00;
14'h175d:data=8'h00;
14'h175e:data=8'h00;
14'h175f:data=8'h00;
14'h1760:data=8'h00;
14'h1761:data=8'h00;
14'h1762:data=8'h00;
14'h1763:data=8'h00;
14'h1764:data=8'h00;
14'h1765:data=8'h00;
14'h1766:data=8'h00;
14'h1767:data=8'h00;
14'h1780:data=8'h00;
14'h1781:data=8'h00;
14'h1782:data=8'h00;
14'h1783:data=8'h00;
14'h1784:data=8'h00;
14'h1785:data=8'h00;
14'h1786:data=8'h00;
14'h1787:data=8'h00;
14'h1788:data=8'h00;
14'h1789:data=8'h00;
14'h178a:data=8'h07;
14'h178b:data=8'hFF;
14'h178c:data=8'hF8;
14'h178d:data=8'h00;
14'h178e:data=8'h00;
14'h178f:data=8'h00;
14'h1790:data=8'h00;
14'h1791:data=8'h07;
14'h1792:data=8'hFF;
14'h1793:data=8'hFE;
14'h1794:data=8'h00;
14'h1795:data=8'h00;
14'h1796:data=8'h00;
14'h1797:data=8'h00;
14'h1798:data=8'h00;
14'h1799:data=8'h00;
14'h179a:data=8'h00;
14'h179b:data=8'h00;
14'h179c:data=8'h00;
14'h179d:data=8'h00;
14'h179e:data=8'h00;
14'h179f:data=8'h00;
14'h17a0:data=8'h00;
14'h17a1:data=8'h00;
14'h17a2:data=8'h00;
14'h17a3:data=8'h00;
14'h17a4:data=8'h00;
14'h17a5:data=8'h00;
14'h17a6:data=8'h00;
14'h17a7:data=8'h00;
14'h17c0:data=8'h00;
14'h17c1:data=8'h0F;
14'h17c2:data=8'hFF;
14'h17c3:data=8'hFC;
14'h17c4:data=8'h00;
14'h17c5:data=8'h00;
14'h17c6:data=8'h00;
14'h17c7:data=8'h00;
14'h17c8:data=8'h00;
14'h17c9:data=8'h00;
14'h17ca:data=8'h07;
14'h17cb:data=8'hFF;
14'h17cc:data=8'hF8;
14'h17cd:data=8'h00;
14'h17ce:data=8'h00;
14'h17cf:data=8'h00;
14'h17d0:data=8'h00;
14'h17d1:data=8'h07;
14'h17d2:data=8'hFF;
14'h17d3:data=8'hFE;
14'h17d4:data=8'h00;
14'h17d5:data=8'h00;
14'h17d6:data=8'h00;
14'h17d7:data=8'h00;
14'h17d8:data=8'h00;
14'h17d9:data=8'h1F;
14'h17da:data=8'hFF;
14'h17db:data=8'hFF;
14'h17dc:data=8'hF8;
14'h17dd:data=8'h00;
14'h17de:data=8'h00;
14'h17df:data=8'h00;
14'h17e0:data=8'h00;
14'h17e1:data=8'h00;
14'h17e2:data=8'h7F;
14'h17e3:data=8'hFF;
14'h17e4:data=8'hFF;
14'h17e5:data=8'hFC;
14'h17e6:data=8'h00;
14'h17e7:data=8'h00;
14'h1800:data=8'h00;
14'h1801:data=8'h0F;
14'h1802:data=8'hFF;
14'h1803:data=8'hFC;
14'h1804:data=8'h00;
14'h1805:data=8'h00;
14'h1806:data=8'h00;
14'h1807:data=8'h00;
14'h1808:data=8'h00;
14'h1809:data=8'h00;
14'h180a:data=8'h07;
14'h180b:data=8'hFF;
14'h180c:data=8'hF8;
14'h180d:data=8'h00;
14'h180e:data=8'h00;
14'h180f:data=8'h00;
14'h1810:data=8'h00;
14'h1811:data=8'h07;
14'h1812:data=8'hFF;
14'h1813:data=8'hFE;
14'h1814:data=8'h00;
14'h1815:data=8'h00;
14'h1816:data=8'h00;
14'h1817:data=8'h00;
14'h1818:data=8'h00;
14'h1819:data=8'h1F;
14'h181a:data=8'hFF;
14'h181b:data=8'hFF;
14'h181c:data=8'hF8;
14'h181d:data=8'h00;
14'h181e:data=8'h00;
14'h181f:data=8'h00;
14'h1820:data=8'h00;
14'h1821:data=8'h00;
14'h1822:data=8'h7F;
14'h1823:data=8'hFF;
14'h1824:data=8'hFF;
14'h1825:data=8'hFC;
14'h1826:data=8'h00;
14'h1827:data=8'h00;
14'h1840:data=8'h00;
14'h1841:data=8'h0F;
14'h1842:data=8'hFF;
14'h1843:data=8'hFC;
14'h1844:data=8'h00;
14'h1845:data=8'h00;
14'h1846:data=8'h00;
14'h1847:data=8'h00;
14'h1848:data=8'h00;
14'h1849:data=8'h3F;
14'h184a:data=8'hFF;
14'h184b:data=8'hFF;
14'h184c:data=8'hF8;
14'h184d:data=8'h00;
14'h184e:data=8'h00;
14'h184f:data=8'h00;
14'h1850:data=8'h00;
14'h1851:data=8'h07;
14'h1852:data=8'hFF;
14'h1853:data=8'hFE;
14'h1854:data=8'h00;
14'h1855:data=8'h00;
14'h1856:data=8'h00;
14'h1857:data=8'h00;
14'h1858:data=8'h00;
14'h1859:data=8'h1F;
14'h185a:data=8'hFF;
14'h185b:data=8'hFF;
14'h185c:data=8'hF8;
14'h185d:data=8'h00;
14'h185e:data=8'h00;
14'h185f:data=8'h00;
14'h1860:data=8'h00;
14'h1861:data=8'h00;
14'h1862:data=8'h7F;
14'h1863:data=8'hFF;
14'h1864:data=8'hFF;
14'h1865:data=8'hFC;
14'h1866:data=8'h00;
14'h1867:data=8'h00;
14'h1880:data=8'h00;
14'h1881:data=8'h0F;
14'h1882:data=8'hFF;
14'h1883:data=8'hFC;
14'h1884:data=8'h00;
14'h1885:data=8'h00;
14'h1886:data=8'h00;
14'h1887:data=8'h00;
14'h1888:data=8'h00;
14'h1889:data=8'h3F;
14'h188a:data=8'hFF;
14'h188b:data=8'hFF;
14'h188c:data=8'hF8;
14'h188d:data=8'h00;
14'h188e:data=8'h00;
14'h188f:data=8'h00;
14'h1890:data=8'h00;
14'h1891:data=8'h07;
14'h1892:data=8'hFF;
14'h1893:data=8'hFF;
14'h1894:data=8'hF8;
14'h1895:data=8'h00;
14'h1896:data=8'h00;
14'h1897:data=8'h00;
14'h1898:data=8'h00;
14'h1899:data=8'h1F;
14'h189a:data=8'hFF;
14'h189b:data=8'hFF;
14'h189c:data=8'hF8;
14'h189d:data=8'h00;
14'h189e:data=8'h00;
14'h189f:data=8'h00;
14'h18a0:data=8'h00;
14'h18a1:data=8'h00;
14'h18a2:data=8'h7F;
14'h18a3:data=8'hFF;
14'h18a4:data=8'hFF;
14'h18a5:data=8'hFC;
14'h18a6:data=8'h00;
14'h18a7:data=8'h00;
14'h18c0:data=8'h00;
14'h18c1:data=8'h0F;
14'h18c2:data=8'hFF;
14'h18c3:data=8'hFC;
14'h18c4:data=8'h00;
14'h18c5:data=8'h00;
14'h18c6:data=8'h00;
14'h18c7:data=8'h00;
14'h18c8:data=8'h00;
14'h18c9:data=8'h3F;
14'h18ca:data=8'hFF;
14'h18cb:data=8'hFF;
14'h18cc:data=8'hF8;
14'h18cd:data=8'h00;
14'h18ce:data=8'h00;
14'h18cf:data=8'h00;
14'h18d0:data=8'h00;
14'h18d1:data=8'h07;
14'h18d2:data=8'hFF;
14'h18d3:data=8'hFF;
14'h18d4:data=8'hF8;
14'h18d5:data=8'h00;
14'h18d6:data=8'h00;
14'h18d7:data=8'h00;
14'h18d8:data=8'h00;
14'h18d9:data=8'h1F;
14'h18da:data=8'hFF;
14'h18db:data=8'hFF;
14'h18dc:data=8'hF8;
14'h18dd:data=8'h00;
14'h18de:data=8'h00;
14'h18df:data=8'h00;
14'h18e0:data=8'h00;
14'h18e1:data=8'h00;
14'h18e2:data=8'h7F;
14'h18e3:data=8'hFF;
14'h18e4:data=8'hFF;
14'h18e5:data=8'hFC;
14'h18e6:data=8'h00;
14'h18e7:data=8'h00;
14'h1900:data=8'h00;
14'h1901:data=8'h0F;
14'h1902:data=8'hFF;
14'h1903:data=8'hFC;
14'h1904:data=8'h00;
14'h1905:data=8'h00;
14'h1906:data=8'h00;
14'h1907:data=8'h00;
14'h1908:data=8'h00;
14'h1909:data=8'h3F;
14'h190a:data=8'hFF;
14'h190b:data=8'hFF;
14'h190c:data=8'hF8;
14'h190d:data=8'h00;
14'h190e:data=8'h00;
14'h190f:data=8'h00;
14'h1910:data=8'h00;
14'h1911:data=8'h07;
14'h1912:data=8'hFF;
14'h1913:data=8'hFF;
14'h1914:data=8'hF8;
14'h1915:data=8'h00;
14'h1916:data=8'h00;
14'h1917:data=8'h00;
14'h1918:data=8'h00;
14'h1919:data=8'h1F;
14'h191a:data=8'hFF;
14'h191b:data=8'hFF;
14'h191c:data=8'hF8;
14'h191d:data=8'h00;
14'h191e:data=8'h00;
14'h191f:data=8'h00;
14'h1920:data=8'h00;
14'h1921:data=8'h00;
14'h1922:data=8'h7F;
14'h1923:data=8'hFF;
14'h1924:data=8'hFF;
14'h1925:data=8'hFC;
14'h1926:data=8'h00;
14'h1927:data=8'h00;
14'h1940:data=8'h00;
14'h1941:data=8'h07;
14'h1942:data=8'hFF;
14'h1943:data=8'hFC;
14'h1944:data=8'h00;
14'h1945:data=8'h00;
14'h1946:data=8'h00;
14'h1947:data=8'h00;
14'h1948:data=8'h00;
14'h1949:data=8'h3F;
14'h194a:data=8'hFF;
14'h194b:data=8'hFF;
14'h194c:data=8'hF8;
14'h194d:data=8'h00;
14'h194e:data=8'h00;
14'h194f:data=8'h00;
14'h1950:data=8'h00;
14'h1951:data=8'h07;
14'h1952:data=8'hFF;
14'h1953:data=8'hFF;
14'h1954:data=8'hF8;
14'h1955:data=8'h00;
14'h1956:data=8'h00;
14'h1957:data=8'h00;
14'h1958:data=8'h00;
14'h1959:data=8'h1F;
14'h195a:data=8'hFF;
14'h195b:data=8'hFF;
14'h195c:data=8'hF8;
14'h195d:data=8'h00;
14'h195e:data=8'h00;
14'h195f:data=8'h00;
14'h1960:data=8'h00;
14'h1961:data=8'h00;
14'h1962:data=8'h7F;
14'h1963:data=8'hFF;
14'h1964:data=8'hFF;
14'h1965:data=8'hFC;
14'h1966:data=8'h00;
14'h1967:data=8'h00;
14'h1980:data=8'h00;
14'h1981:data=8'h07;
14'h1982:data=8'hFF;
14'h1983:data=8'hFC;
14'h1984:data=8'h00;
14'h1985:data=8'h00;
14'h1986:data=8'h00;
14'h1987:data=8'h00;
14'h1988:data=8'h00;
14'h1989:data=8'h3F;
14'h198a:data=8'hFF;
14'h198b:data=8'hFF;
14'h198c:data=8'hF8;
14'h198d:data=8'h00;
14'h198e:data=8'h00;
14'h198f:data=8'h00;
14'h1990:data=8'h00;
14'h1991:data=8'h07;
14'h1992:data=8'hFF;
14'h1993:data=8'hFF;
14'h1994:data=8'hF8;
14'h1995:data=8'h00;
14'h1996:data=8'h00;
14'h1997:data=8'h00;
14'h1998:data=8'h00;
14'h1999:data=8'h1F;
14'h199a:data=8'hFF;
14'h199b:data=8'hFF;
14'h199c:data=8'hF8;
14'h199d:data=8'h00;
14'h199e:data=8'h00;
14'h199f:data=8'h00;
14'h19a0:data=8'h00;
14'h19a1:data=8'h00;
14'h19a2:data=8'h7F;
14'h19a3:data=8'hFF;
14'h19a4:data=8'hFF;
14'h19a5:data=8'hFC;
14'h19a6:data=8'h00;
14'h19a7:data=8'h00;
14'h19c0:data=8'h00;
14'h19c1:data=8'h07;
14'h19c2:data=8'hFF;
14'h19c3:data=8'hFC;
14'h19c4:data=8'h00;
14'h19c5:data=8'h00;
14'h19c6:data=8'h00;
14'h19c7:data=8'h00;
14'h19c8:data=8'h00;
14'h19c9:data=8'h3F;
14'h19ca:data=8'hFF;
14'h19cb:data=8'hFF;
14'h19cc:data=8'hF8;
14'h19cd:data=8'h00;
14'h19ce:data=8'h00;
14'h19cf:data=8'h00;
14'h19d0:data=8'h00;
14'h19d1:data=8'h07;
14'h19d2:data=8'hFF;
14'h19d3:data=8'hFF;
14'h19d4:data=8'hFC;
14'h19d5:data=8'h00;
14'h19d6:data=8'h00;
14'h19d7:data=8'h00;
14'h19d8:data=8'h00;
14'h19d9:data=8'h1F;
14'h19da:data=8'hFF;
14'h19db:data=8'hFF;
14'h19dc:data=8'hF8;
14'h19dd:data=8'h00;
14'h19de:data=8'h00;
14'h19df:data=8'h00;
14'h19e0:data=8'h00;
14'h19e1:data=8'h00;
14'h19e2:data=8'h7F;
14'h19e3:data=8'hFF;
14'h19e4:data=8'hFF;
14'h19e5:data=8'hFC;
14'h19e6:data=8'h00;
14'h19e7:data=8'h00;
14'h1a00:data=8'h00;
14'h1a01:data=8'h07;
14'h1a02:data=8'hFF;
14'h1a03:data=8'hFC;
14'h1a04:data=8'h00;
14'h1a05:data=8'h00;
14'h1a06:data=8'h00;
14'h1a07:data=8'h00;
14'h1a08:data=8'h00;
14'h1a09:data=8'h3F;
14'h1a0a:data=8'hFF;
14'h1a0b:data=8'hFF;
14'h1a0c:data=8'hF8;
14'h1a0d:data=8'h00;
14'h1a0e:data=8'h00;
14'h1a0f:data=8'h00;
14'h1a10:data=8'h00;
14'h1a11:data=8'h07;
14'h1a12:data=8'hFF;
14'h1a13:data=8'hFF;
14'h1a14:data=8'hFC;
14'h1a15:data=8'h00;
14'h1a16:data=8'h00;
14'h1a17:data=8'h00;
14'h1a18:data=8'h00;
14'h1a19:data=8'h1F;
14'h1a1a:data=8'hFF;
14'h1a1b:data=8'hFF;
14'h1a1c:data=8'hF8;
14'h1a1d:data=8'h00;
14'h1a1e:data=8'h00;
14'h1a1f:data=8'h00;
14'h1a20:data=8'h00;
14'h1a21:data=8'h00;
14'h1a22:data=8'h3F;
14'h1a23:data=8'hFF;
14'h1a24:data=8'hFF;
14'h1a25:data=8'hFC;
14'h1a26:data=8'h00;
14'h1a27:data=8'h00;
14'h1a40:data=8'h00;
14'h1a41:data=8'h07;
14'h1a42:data=8'hFF;
14'h1a43:data=8'hFC;
14'h1a44:data=8'h00;
14'h1a45:data=8'h00;
14'h1a46:data=8'h00;
14'h1a47:data=8'h00;
14'h1a48:data=8'h00;
14'h1a49:data=8'h3F;
14'h1a4a:data=8'hFF;
14'h1a4b:data=8'hFF;
14'h1a4c:data=8'hF8;
14'h1a4d:data=8'h00;
14'h1a4e:data=8'h00;
14'h1a4f:data=8'h00;
14'h1a50:data=8'h00;
14'h1a51:data=8'h07;
14'h1a52:data=8'hFF;
14'h1a53:data=8'hFF;
14'h1a54:data=8'hFC;
14'h1a55:data=8'h00;
14'h1a56:data=8'h00;
14'h1a57:data=8'h00;
14'h1a58:data=8'h00;
14'h1a59:data=8'h1F;
14'h1a5a:data=8'hFF;
14'h1a5b:data=8'hFF;
14'h1a5c:data=8'hF8;
14'h1a5d:data=8'h00;
14'h1a5e:data=8'h00;
14'h1a5f:data=8'h00;
14'h1a60:data=8'h00;
14'h1a61:data=8'h00;
14'h1a62:data=8'h3F;
14'h1a63:data=8'hFF;
14'h1a64:data=8'hFF;
14'h1a65:data=8'hFC;
14'h1a66:data=8'h00;
14'h1a67:data=8'h00;
14'h1a80:data=8'h00;
14'h1a81:data=8'h07;
14'h1a82:data=8'hFF;
14'h1a83:data=8'hFC;
14'h1a84:data=8'h00;
14'h1a85:data=8'h00;
14'h1a86:data=8'h00;
14'h1a87:data=8'h00;
14'h1a88:data=8'h00;
14'h1a89:data=8'h3F;
14'h1a8a:data=8'hFF;
14'h1a8b:data=8'hFF;
14'h1a8c:data=8'hF8;
14'h1a8d:data=8'h00;
14'h1a8e:data=8'h00;
14'h1a8f:data=8'h00;
14'h1a90:data=8'h00;
14'h1a91:data=8'h07;
14'h1a92:data=8'hFF;
14'h1a93:data=8'hFF;
14'h1a94:data=8'hFC;
14'h1a95:data=8'h00;
14'h1a96:data=8'h00;
14'h1a97:data=8'h00;
14'h1a98:data=8'h00;
14'h1a99:data=8'h1F;
14'h1a9a:data=8'hFF;
14'h1a9b:data=8'hFF;
14'h1a9c:data=8'hF8;
14'h1a9d:data=8'h00;
14'h1a9e:data=8'h00;
14'h1a9f:data=8'h00;
14'h1aa0:data=8'h00;
14'h1aa1:data=8'h00;
14'h1aa2:data=8'h3F;
14'h1aa3:data=8'hFF;
14'h1aa4:data=8'hFF;
14'h1aa5:data=8'hFC;
14'h1aa6:data=8'h00;
14'h1aa7:data=8'h00;
14'h1ac0:data=8'h00;
14'h1ac1:data=8'h07;
14'h1ac2:data=8'hFF;
14'h1ac3:data=8'hFC;
14'h1ac4:data=8'h00;
14'h1ac5:data=8'h00;
14'h1ac6:data=8'h00;
14'h1ac7:data=8'h00;
14'h1ac8:data=8'h00;
14'h1ac9:data=8'h3F;
14'h1aca:data=8'hFF;
14'h1acb:data=8'hFF;
14'h1acc:data=8'hF8;
14'h1acd:data=8'h00;
14'h1ace:data=8'h00;
14'h1acf:data=8'h00;
14'h1ad0:data=8'h00;
14'h1ad1:data=8'h07;
14'h1ad2:data=8'hFF;
14'h1ad3:data=8'hFF;
14'h1ad4:data=8'hFC;
14'h1ad5:data=8'h00;
14'h1ad6:data=8'h00;
14'h1ad7:data=8'h00;
14'h1ad8:data=8'h00;
14'h1ad9:data=8'h1F;
14'h1ada:data=8'hFF;
14'h1adb:data=8'hFF;
14'h1adc:data=8'hF8;
14'h1add:data=8'h00;
14'h1ade:data=8'h00;
14'h1adf:data=8'h00;
14'h1ae0:data=8'h00;
14'h1ae1:data=8'h00;
14'h1ae2:data=8'h3F;
14'h1ae3:data=8'hFF;
14'h1ae4:data=8'hFF;
14'h1ae5:data=8'hFC;
14'h1ae6:data=8'h00;
14'h1ae7:data=8'h00;
14'h1b00:data=8'h00;
14'h1b01:data=8'h07;
14'h1b02:data=8'hFF;
14'h1b03:data=8'hFE;
14'h1b04:data=8'h00;
14'h1b05:data=8'h00;
14'h1b06:data=8'h00;
14'h1b07:data=8'h00;
14'h1b08:data=8'h00;
14'h1b09:data=8'h3F;
14'h1b0a:data=8'hFF;
14'h1b0b:data=8'hFF;
14'h1b0c:data=8'hF8;
14'h1b0d:data=8'h00;
14'h1b0e:data=8'h00;
14'h1b0f:data=8'h00;
14'h1b10:data=8'h00;
14'h1b11:data=8'h07;
14'h1b12:data=8'hFF;
14'h1b13:data=8'hFF;
14'h1b14:data=8'hFC;
14'h1b15:data=8'h00;
14'h1b16:data=8'h00;
14'h1b17:data=8'h00;
14'h1b18:data=8'h00;
14'h1b19:data=8'h1F;
14'h1b1a:data=8'hFF;
14'h1b1b:data=8'hFF;
14'h1b1c:data=8'hF8;
14'h1b1d:data=8'h00;
14'h1b1e:data=8'h00;
14'h1b1f:data=8'h00;
14'h1b20:data=8'h00;
14'h1b21:data=8'h00;
14'h1b22:data=8'h3F;
14'h1b23:data=8'hFF;
14'h1b24:data=8'hFF;
14'h1b25:data=8'hFC;
14'h1b26:data=8'h00;
14'h1b27:data=8'h00;
14'h1b40:data=8'h00;
14'h1b41:data=8'h07;
14'h1b42:data=8'hFF;
14'h1b43:data=8'hFE;
14'h1b44:data=8'h00;
14'h1b45:data=8'h00;
14'h1b46:data=8'h00;
14'h1b47:data=8'h00;
14'h1b48:data=8'h00;
14'h1b49:data=8'h3F;
14'h1b4a:data=8'hFF;
14'h1b4b:data=8'hFF;
14'h1b4c:data=8'hF8;
14'h1b4d:data=8'h00;
14'h1b4e:data=8'h00;
14'h1b4f:data=8'h00;
14'h1b50:data=8'h00;
14'h1b51:data=8'h07;
14'h1b52:data=8'hFF;
14'h1b53:data=8'hFF;
14'h1b54:data=8'hFC;
14'h1b55:data=8'h00;
14'h1b56:data=8'h00;
14'h1b57:data=8'h00;
14'h1b58:data=8'h00;
14'h1b59:data=8'h1F;
14'h1b5a:data=8'hFF;
14'h1b5b:data=8'hFF;
14'h1b5c:data=8'hF8;
14'h1b5d:data=8'h00;
14'h1b5e:data=8'h00;
14'h1b5f:data=8'h00;
14'h1b60:data=8'h00;
14'h1b61:data=8'h00;
14'h1b62:data=8'h3F;
14'h1b63:data=8'hFF;
14'h1b64:data=8'hFF;
14'h1b65:data=8'hFC;
14'h1b66:data=8'h00;
14'h1b67:data=8'h00;
14'h1b80:data=8'h00;
14'h1b81:data=8'h07;
14'h1b82:data=8'hFF;
14'h1b83:data=8'hFE;
14'h1b84:data=8'h00;
14'h1b85:data=8'h00;
14'h1b86:data=8'h00;
14'h1b87:data=8'h00;
14'h1b88:data=8'h00;
14'h1b89:data=8'h3F;
14'h1b8a:data=8'hFF;
14'h1b8b:data=8'hFF;
14'h1b8c:data=8'hF8;
14'h1b8d:data=8'h00;
14'h1b8e:data=8'h00;
14'h1b8f:data=8'h00;
14'h1b90:data=8'h00;
14'h1b91:data=8'h07;
14'h1b92:data=8'hFF;
14'h1b93:data=8'hFF;
14'h1b94:data=8'hFC;
14'h1b95:data=8'h00;
14'h1b96:data=8'h00;
14'h1b97:data=8'h00;
14'h1b98:data=8'h00;
14'h1b99:data=8'h1F;
14'h1b9a:data=8'hFF;
14'h1b9b:data=8'hFF;
14'h1b9c:data=8'hF8;
14'h1b9d:data=8'h00;
14'h1b9e:data=8'h00;
14'h1b9f:data=8'h00;
14'h1ba0:data=8'h00;
14'h1ba1:data=8'h00;
14'h1ba2:data=8'h3F;
14'h1ba3:data=8'hFF;
14'h1ba4:data=8'hFF;
14'h1ba5:data=8'hFC;
14'h1ba6:data=8'h00;
14'h1ba7:data=8'h00;
14'h1bc0:data=8'h00;
14'h1bc1:data=8'h07;
14'h1bc2:data=8'hFF;
14'h1bc3:data=8'hFE;
14'h1bc4:data=8'h00;
14'h1bc5:data=8'h00;
14'h1bc6:data=8'h00;
14'h1bc7:data=8'h00;
14'h1bc8:data=8'h00;
14'h1bc9:data=8'h3F;
14'h1bca:data=8'hFF;
14'h1bcb:data=8'hFF;
14'h1bcc:data=8'hF8;
14'h1bcd:data=8'h00;
14'h1bce:data=8'h00;
14'h1bcf:data=8'h00;
14'h1bd0:data=8'h00;
14'h1bd1:data=8'h07;
14'h1bd2:data=8'hFF;
14'h1bd3:data=8'hFF;
14'h1bd4:data=8'hFC;
14'h1bd5:data=8'h00;
14'h1bd6:data=8'h00;
14'h1bd7:data=8'h00;
14'h1bd8:data=8'h00;
14'h1bd9:data=8'h1F;
14'h1bda:data=8'hFF;
14'h1bdb:data=8'hFF;
14'h1bdc:data=8'hF8;
14'h1bdd:data=8'h00;
14'h1bde:data=8'h00;
14'h1bdf:data=8'h00;
14'h1be0:data=8'h00;
14'h1be1:data=8'h00;
14'h1be2:data=8'h3F;
14'h1be3:data=8'hFF;
14'h1be4:data=8'hFF;
14'h1be5:data=8'hFC;
14'h1be6:data=8'h00;
14'h1be7:data=8'h00;
14'h1c00:data=8'h00;
14'h1c01:data=8'h07;
14'h1c02:data=8'hFF;
14'h1c03:data=8'hFE;
14'h1c04:data=8'h00;
14'h1c05:data=8'h00;
14'h1c06:data=8'h00;
14'h1c07:data=8'h00;
14'h1c08:data=8'h00;
14'h1c09:data=8'h3F;
14'h1c0a:data=8'hFF;
14'h1c0b:data=8'hFF;
14'h1c0c:data=8'hF8;
14'h1c0d:data=8'h00;
14'h1c0e:data=8'h00;
14'h1c0f:data=8'h00;
14'h1c10:data=8'h00;
14'h1c11:data=8'h07;
14'h1c12:data=8'hFF;
14'h1c13:data=8'hFF;
14'h1c14:data=8'hFC;
14'h1c15:data=8'h00;
14'h1c16:data=8'h00;
14'h1c17:data=8'h00;
14'h1c18:data=8'h00;
14'h1c19:data=8'h1F;
14'h1c1a:data=8'hFF;
14'h1c1b:data=8'hFF;
14'h1c1c:data=8'hF8;
14'h1c1d:data=8'h00;
14'h1c1e:data=8'h00;
14'h1c1f:data=8'h00;
14'h1c20:data=8'h00;
14'h1c21:data=8'h00;
14'h1c22:data=8'h3F;
14'h1c23:data=8'hFF;
14'h1c24:data=8'hFF;
14'h1c25:data=8'hFC;
14'h1c26:data=8'h00;
14'h1c27:data=8'h00;
14'h1c40:data=8'h00;
14'h1c41:data=8'h07;
14'h1c42:data=8'hFF;
14'h1c43:data=8'hFE;
14'h1c44:data=8'h00;
14'h1c45:data=8'h00;
14'h1c46:data=8'h00;
14'h1c47:data=8'h00;
14'h1c48:data=8'h00;
14'h1c49:data=8'h3F;
14'h1c4a:data=8'hFF;
14'h1c4b:data=8'hFF;
14'h1c4c:data=8'hF8;
14'h1c4d:data=8'h00;
14'h1c4e:data=8'h00;
14'h1c4f:data=8'h00;
14'h1c50:data=8'h00;
14'h1c51:data=8'h07;
14'h1c52:data=8'hFF;
14'h1c53:data=8'hFF;
14'h1c54:data=8'hFC;
14'h1c55:data=8'h00;
14'h1c56:data=8'h00;
14'h1c57:data=8'h00;
14'h1c58:data=8'h00;
14'h1c59:data=8'h1F;
14'h1c5a:data=8'hFF;
14'h1c5b:data=8'hFF;
14'h1c5c:data=8'hF8;
14'h1c5d:data=8'h00;
14'h1c5e:data=8'h00;
14'h1c5f:data=8'h00;
14'h1c60:data=8'h00;
14'h1c61:data=8'h00;
14'h1c62:data=8'h3F;
14'h1c63:data=8'hFF;
14'h1c64:data=8'hFF;
14'h1c65:data=8'hFC;
14'h1c66:data=8'h00;
14'h1c67:data=8'h00;
14'h1c80:data=8'h00;
14'h1c81:data=8'h07;
14'h1c82:data=8'hFF;
14'h1c83:data=8'hFE;
14'h1c84:data=8'h00;
14'h1c85:data=8'h00;
14'h1c86:data=8'h00;
14'h1c87:data=8'h00;
14'h1c88:data=8'h00;
14'h1c89:data=8'h1F;
14'h1c8a:data=8'hFF;
14'h1c8b:data=8'hFF;
14'h1c8c:data=8'hF8;
14'h1c8d:data=8'h00;
14'h1c8e:data=8'h00;
14'h1c8f:data=8'h00;
14'h1c90:data=8'h00;
14'h1c91:data=8'h07;
14'h1c92:data=8'hFF;
14'h1c93:data=8'hFF;
14'h1c94:data=8'hFC;
14'h1c95:data=8'h00;
14'h1c96:data=8'h00;
14'h1c97:data=8'h00;
14'h1c98:data=8'h00;
14'h1c99:data=8'h1F;
14'h1c9a:data=8'hFF;
14'h1c9b:data=8'hFF;
14'h1c9c:data=8'hF8;
14'h1c9d:data=8'h00;
14'h1c9e:data=8'h00;
14'h1c9f:data=8'h00;
14'h1ca0:data=8'h00;
14'h1ca1:data=8'h00;
14'h1ca2:data=8'h3F;
14'h1ca3:data=8'hFF;
14'h1ca4:data=8'hFF;
14'h1ca5:data=8'hFC;
14'h1ca6:data=8'h00;
14'h1ca7:data=8'h00;
14'h1cc0:data=8'h00;
14'h1cc1:data=8'h07;
14'h1cc2:data=8'hFF;
14'h1cc3:data=8'hFE;
14'h1cc4:data=8'h00;
14'h1cc5:data=8'h00;
14'h1cc6:data=8'h00;
14'h1cc7:data=8'h00;
14'h1cc8:data=8'h00;
14'h1cc9:data=8'h1F;
14'h1cca:data=8'hFF;
14'h1ccb:data=8'hFF;
14'h1ccc:data=8'hF8;
14'h1ccd:data=8'h00;
14'h1cce:data=8'h00;
14'h1ccf:data=8'h00;
14'h1cd0:data=8'h00;
14'h1cd1:data=8'h07;
14'h1cd2:data=8'hFF;
14'h1cd3:data=8'hFF;
14'h1cd4:data=8'hFC;
14'h1cd5:data=8'h00;
14'h1cd6:data=8'h00;
14'h1cd7:data=8'h00;
14'h1cd8:data=8'h00;
14'h1cd9:data=8'h1F;
14'h1cda:data=8'hFF;
14'h1cdb:data=8'hFF;
14'h1cdc:data=8'hF8;
14'h1cdd:data=8'h00;
14'h1cde:data=8'h00;
14'h1cdf:data=8'h00;
14'h1ce0:data=8'h00;
14'h1ce1:data=8'h00;
14'h1ce2:data=8'h3F;
14'h1ce3:data=8'hFF;
14'h1ce4:data=8'hFF;
14'h1ce5:data=8'hFC;
14'h1ce6:data=8'h00;
14'h1ce7:data=8'h00;
14'h1d00:data=8'h00;
14'h1d01:data=8'h07;
14'h1d02:data=8'hFF;
14'h1d03:data=8'hFE;
14'h1d04:data=8'h00;
14'h1d05:data=8'h00;
14'h1d06:data=8'h00;
14'h1d07:data=8'h00;
14'h1d08:data=8'h00;
14'h1d09:data=8'h1F;
14'h1d0a:data=8'hFF;
14'h1d0b:data=8'hFF;
14'h1d0c:data=8'hF8;
14'h1d0d:data=8'h00;
14'h1d0e:data=8'h00;
14'h1d0f:data=8'h00;
14'h1d10:data=8'h00;
14'h1d11:data=8'h07;
14'h1d12:data=8'hFF;
14'h1d13:data=8'hFF;
14'h1d14:data=8'hFC;
14'h1d15:data=8'h00;
14'h1d16:data=8'h00;
14'h1d17:data=8'h00;
14'h1d18:data=8'h00;
14'h1d19:data=8'h1F;
14'h1d1a:data=8'hFF;
14'h1d1b:data=8'hFF;
14'h1d1c:data=8'hF8;
14'h1d1d:data=8'h00;
14'h1d1e:data=8'h00;
14'h1d1f:data=8'h00;
14'h1d20:data=8'h00;
14'h1d21:data=8'h00;
14'h1d22:data=8'h3F;
14'h1d23:data=8'hFF;
14'h1d24:data=8'hFF;
14'h1d25:data=8'hFC;
14'h1d26:data=8'h00;
14'h1d27:data=8'h00;
14'h1d40:data=8'h00;
14'h1d41:data=8'h07;
14'h1d42:data=8'hFF;
14'h1d43:data=8'hFE;
14'h1d44:data=8'h00;
14'h1d45:data=8'h00;
14'h1d46:data=8'h00;
14'h1d47:data=8'h00;
14'h1d48:data=8'h00;
14'h1d49:data=8'h1F;
14'h1d4a:data=8'hFF;
14'h1d4b:data=8'hFF;
14'h1d4c:data=8'hF8;
14'h1d4d:data=8'h00;
14'h1d4e:data=8'h00;
14'h1d4f:data=8'h00;
14'h1d50:data=8'h00;
14'h1d51:data=8'h07;
14'h1d52:data=8'hFF;
14'h1d53:data=8'hFF;
14'h1d54:data=8'hFC;
14'h1d55:data=8'h00;
14'h1d56:data=8'h00;
14'h1d57:data=8'h00;
14'h1d58:data=8'h00;
14'h1d59:data=8'h1F;
14'h1d5a:data=8'hFF;
14'h1d5b:data=8'hFF;
14'h1d5c:data=8'hF8;
14'h1d5d:data=8'h00;
14'h1d5e:data=8'h00;
14'h1d5f:data=8'h00;
14'h1d60:data=8'h00;
14'h1d61:data=8'h00;
14'h1d62:data=8'h3F;
14'h1d63:data=8'hFF;
14'h1d64:data=8'hFF;
14'h1d65:data=8'hFC;
14'h1d66:data=8'h00;
14'h1d67:data=8'h00;
14'h1d80:data=8'h00;
14'h1d81:data=8'h07;
14'h1d82:data=8'hFF;
14'h1d83:data=8'hFE;
14'h1d84:data=8'h00;
14'h1d85:data=8'h00;
14'h1d86:data=8'h00;
14'h1d87:data=8'h00;
14'h1d88:data=8'h00;
14'h1d89:data=8'h1F;
14'h1d8a:data=8'hFF;
14'h1d8b:data=8'hFF;
14'h1d8c:data=8'hF8;
14'h1d8d:data=8'h00;
14'h1d8e:data=8'h00;
14'h1d8f:data=8'h00;
14'h1d90:data=8'h00;
14'h1d91:data=8'h07;
14'h1d92:data=8'hFF;
14'h1d93:data=8'hFF;
14'h1d94:data=8'hFC;
14'h1d95:data=8'h00;
14'h1d96:data=8'h00;
14'h1d97:data=8'h00;
14'h1d98:data=8'h00;
14'h1d99:data=8'h1F;
14'h1d9a:data=8'hFF;
14'h1d9b:data=8'hFF;
14'h1d9c:data=8'hF8;
14'h1d9d:data=8'h00;
14'h1d9e:data=8'h00;
14'h1d9f:data=8'h00;
14'h1da0:data=8'h00;
14'h1da1:data=8'h00;
14'h1da2:data=8'h3F;
14'h1da3:data=8'hFF;
14'h1da4:data=8'hFF;
14'h1da5:data=8'hFC;
14'h1da6:data=8'h00;
14'h1da7:data=8'h00;
14'h1dc0:data=8'h00;
14'h1dc1:data=8'h07;
14'h1dc2:data=8'hFF;
14'h1dc3:data=8'hFE;
14'h1dc4:data=8'h00;
14'h1dc5:data=8'h00;
14'h1dc6:data=8'h00;
14'h1dc7:data=8'h00;
14'h1dc8:data=8'h00;
14'h1dc9:data=8'h1F;
14'h1dca:data=8'hFF;
14'h1dcb:data=8'hFF;
14'h1dcc:data=8'hF8;
14'h1dcd:data=8'h00;
14'h1dce:data=8'h00;
14'h1dcf:data=8'h00;
14'h1dd0:data=8'h00;
14'h1dd1:data=8'h07;
14'h1dd2:data=8'hFF;
14'h1dd3:data=8'hFF;
14'h1dd4:data=8'hFC;
14'h1dd5:data=8'h00;
14'h1dd6:data=8'h00;
14'h1dd7:data=8'h00;
14'h1dd8:data=8'h00;
14'h1dd9:data=8'h1F;
14'h1dda:data=8'hFF;
14'h1ddb:data=8'hFF;
14'h1ddc:data=8'hF8;
14'h1ddd:data=8'h00;
14'h1dde:data=8'h00;
14'h1ddf:data=8'h00;
14'h1de0:data=8'h00;
14'h1de1:data=8'h00;
14'h1de2:data=8'h3F;
14'h1de3:data=8'hFF;
14'h1de4:data=8'hFF;
14'h1de5:data=8'hFC;
14'h1de6:data=8'h00;
14'h1de7:data=8'h00;
14'h1e00:data=8'h00;
14'h1e01:data=8'h07;
14'h1e02:data=8'hFF;
14'h1e03:data=8'hFE;
14'h1e04:data=8'h00;
14'h1e05:data=8'h00;
14'h1e06:data=8'h00;
14'h1e07:data=8'h00;
14'h1e08:data=8'h00;
14'h1e09:data=8'h1F;
14'h1e0a:data=8'hFF;
14'h1e0b:data=8'hFF;
14'h1e0c:data=8'hF8;
14'h1e0d:data=8'h00;
14'h1e0e:data=8'h00;
14'h1e0f:data=8'h00;
14'h1e10:data=8'h00;
14'h1e11:data=8'h07;
14'h1e12:data=8'hFF;
14'h1e13:data=8'hFF;
14'h1e14:data=8'hFC;
14'h1e15:data=8'h00;
14'h1e16:data=8'h00;
14'h1e17:data=8'h00;
14'h1e18:data=8'h00;
14'h1e19:data=8'h1F;
14'h1e1a:data=8'hFF;
14'h1e1b:data=8'hFF;
14'h1e1c:data=8'hFF;
14'h1e1d:data=8'hFF;
14'h1e1e:data=8'hFF;
14'h1e1f:data=8'hFF;
14'h1e20:data=8'hFF;
14'h1e21:data=8'hFF;
14'h1e22:data=8'hFF;
14'h1e23:data=8'hFF;
14'h1e24:data=8'hFF;
14'h1e25:data=8'hFC;
14'h1e26:data=8'h00;
14'h1e27:data=8'h00;
14'h1e40:data=8'h00;
14'h1e41:data=8'h07;
14'h1e42:data=8'hFF;
14'h1e43:data=8'hFE;
14'h1e44:data=8'h00;
14'h1e45:data=8'h00;
14'h1e46:data=8'h00;
14'h1e47:data=8'h00;
14'h1e48:data=8'h00;
14'h1e49:data=8'h1F;
14'h1e4a:data=8'hFF;
14'h1e4b:data=8'hFF;
14'h1e4c:data=8'hF8;
14'h1e4d:data=8'h00;
14'h1e4e:data=8'h00;
14'h1e4f:data=8'h00;
14'h1e50:data=8'h00;
14'h1e51:data=8'h07;
14'h1e52:data=8'hFF;
14'h1e53:data=8'hFF;
14'h1e54:data=8'hFC;
14'h1e55:data=8'h00;
14'h1e56:data=8'h00;
14'h1e57:data=8'h00;
14'h1e58:data=8'h00;
14'h1e59:data=8'h1F;
14'h1e5a:data=8'hFF;
14'h1e5b:data=8'hFF;
14'h1e5c:data=8'hFF;
14'h1e5d:data=8'hFF;
14'h1e5e:data=8'hFF;
14'h1e5f:data=8'hFF;
14'h1e60:data=8'hFF;
14'h1e61:data=8'hFF;
14'h1e62:data=8'hFF;
14'h1e63:data=8'hFF;
14'h1e64:data=8'hFF;
14'h1e65:data=8'hFC;
14'h1e66:data=8'h00;
14'h1e67:data=8'h00;
14'h1e80:data=8'h00;
14'h1e81:data=8'h07;
14'h1e82:data=8'hFF;
14'h1e83:data=8'hFE;
14'h1e84:data=8'h00;
14'h1e85:data=8'h00;
14'h1e86:data=8'h00;
14'h1e87:data=8'h00;
14'h1e88:data=8'h00;
14'h1e89:data=8'h1F;
14'h1e8a:data=8'hFF;
14'h1e8b:data=8'hFF;
14'h1e8c:data=8'hF8;
14'h1e8d:data=8'h00;
14'h1e8e:data=8'h00;
14'h1e8f:data=8'h00;
14'h1e90:data=8'h00;
14'h1e91:data=8'h07;
14'h1e92:data=8'hFF;
14'h1e93:data=8'hFF;
14'h1e94:data=8'hFC;
14'h1e95:data=8'h00;
14'h1e96:data=8'h00;
14'h1e97:data=8'h00;
14'h1e98:data=8'h00;
14'h1e99:data=8'h1F;
14'h1e9a:data=8'hFF;
14'h1e9b:data=8'hFF;
14'h1e9c:data=8'hFF;
14'h1e9d:data=8'hFF;
14'h1e9e:data=8'hFF;
14'h1e9f:data=8'hFF;
14'h1ea0:data=8'hFF;
14'h1ea1:data=8'hFF;
14'h1ea2:data=8'hFF;
14'h1ea3:data=8'hFF;
14'h1ea4:data=8'hFF;
14'h1ea5:data=8'hFC;
14'h1ea6:data=8'h00;
14'h1ea7:data=8'h00;
14'h1ec0:data=8'h00;
14'h1ec1:data=8'h07;
14'h1ec2:data=8'hFF;
14'h1ec3:data=8'hFE;
14'h1ec4:data=8'h00;
14'h1ec5:data=8'h00;
14'h1ec6:data=8'h00;
14'h1ec7:data=8'h00;
14'h1ec8:data=8'h00;
14'h1ec9:data=8'h1F;
14'h1eca:data=8'hFF;
14'h1ecb:data=8'hFF;
14'h1ecc:data=8'hF8;
14'h1ecd:data=8'h00;
14'h1ece:data=8'h00;
14'h1ecf:data=8'h00;
14'h1ed0:data=8'h00;
14'h1ed1:data=8'h07;
14'h1ed2:data=8'hFF;
14'h1ed3:data=8'hFF;
14'h1ed4:data=8'hFC;
14'h1ed5:data=8'h00;
14'h1ed6:data=8'h00;
14'h1ed7:data=8'h00;
14'h1ed8:data=8'h00;
14'h1ed9:data=8'h1F;
14'h1eda:data=8'hFF;
14'h1edb:data=8'hFF;
14'h1edc:data=8'hFF;
14'h1edd:data=8'hFF;
14'h1ede:data=8'hFF;
14'h1edf:data=8'hFF;
14'h1ee0:data=8'hFF;
14'h1ee1:data=8'hFF;
14'h1ee2:data=8'hFF;
14'h1ee3:data=8'hFF;
14'h1ee4:data=8'hFF;
14'h1ee5:data=8'hFC;
14'h1ee6:data=8'h00;
14'h1ee7:data=8'h00;
14'h1f00:data=8'h00;
14'h1f01:data=8'h03;
14'h1f02:data=8'hFF;
14'h1f03:data=8'hFE;
14'h1f04:data=8'h00;
14'h1f05:data=8'h00;
14'h1f06:data=8'h00;
14'h1f07:data=8'h00;
14'h1f08:data=8'h00;
14'h1f09:data=8'h1F;
14'h1f0a:data=8'hFF;
14'h1f0b:data=8'hFF;
14'h1f0c:data=8'hF8;
14'h1f0d:data=8'h00;
14'h1f0e:data=8'h00;
14'h1f0f:data=8'h00;
14'h1f10:data=8'h00;
14'h1f11:data=8'h07;
14'h1f12:data=8'hFF;
14'h1f13:data=8'hFF;
14'h1f14:data=8'hFC;
14'h1f15:data=8'h00;
14'h1f16:data=8'h00;
14'h1f17:data=8'h00;
14'h1f18:data=8'h00;
14'h1f19:data=8'h1F;
14'h1f1a:data=8'hFF;
14'h1f1b:data=8'hFF;
14'h1f1c:data=8'hFF;
14'h1f1d:data=8'hFF;
14'h1f1e:data=8'hFF;
14'h1f1f:data=8'hFF;
14'h1f20:data=8'hFF;
14'h1f21:data=8'hFF;
14'h1f22:data=8'hFF;
14'h1f23:data=8'hFF;
14'h1f24:data=8'hFF;
14'h1f25:data=8'hFC;
14'h1f26:data=8'h00;
14'h1f27:data=8'h00;
14'h1f40:data=8'h00;
14'h1f41:data=8'h03;
14'h1f42:data=8'hFF;
14'h1f43:data=8'hFE;
14'h1f44:data=8'h00;
14'h1f45:data=8'h00;
14'h1f46:data=8'h00;
14'h1f47:data=8'h00;
14'h1f48:data=8'h00;
14'h1f49:data=8'h1F;
14'h1f4a:data=8'hFF;
14'h1f4b:data=8'hFF;
14'h1f4c:data=8'hF8;
14'h1f4d:data=8'h00;
14'h1f4e:data=8'h00;
14'h1f4f:data=8'h00;
14'h1f50:data=8'h00;
14'h1f51:data=8'h07;
14'h1f52:data=8'hFF;
14'h1f53:data=8'hFF;
14'h1f54:data=8'hFC;
14'h1f55:data=8'h00;
14'h1f56:data=8'h00;
14'h1f57:data=8'h00;
14'h1f58:data=8'h00;
14'h1f59:data=8'h1F;
14'h1f5a:data=8'hFF;
14'h1f5b:data=8'hFF;
14'h1f5c:data=8'hFF;
14'h1f5d:data=8'hFF;
14'h1f5e:data=8'hFF;
14'h1f5f:data=8'hFF;
14'h1f60:data=8'hFF;
14'h1f61:data=8'hFF;
14'h1f62:data=8'hFF;
14'h1f63:data=8'hFF;
14'h1f64:data=8'hFF;
14'h1f65:data=8'hFC;
14'h1f66:data=8'h00;
14'h1f67:data=8'h00;
14'h1f80:data=8'h00;
14'h1f81:data=8'h03;
14'h1f82:data=8'hFF;
14'h1f83:data=8'hFE;
14'h1f84:data=8'h00;
14'h1f85:data=8'h00;
14'h1f86:data=8'h00;
14'h1f87:data=8'h00;
14'h1f88:data=8'h00;
14'h1f89:data=8'h1F;
14'h1f8a:data=8'hFF;
14'h1f8b:data=8'hFF;
14'h1f8c:data=8'hF8;
14'h1f8d:data=8'h00;
14'h1f8e:data=8'h00;
14'h1f8f:data=8'h00;
14'h1f90:data=8'h00;
14'h1f91:data=8'h07;
14'h1f92:data=8'hFF;
14'h1f93:data=8'hFF;
14'h1f94:data=8'hFC;
14'h1f95:data=8'h00;
14'h1f96:data=8'h00;
14'h1f97:data=8'h00;
14'h1f98:data=8'h00;
14'h1f99:data=8'h1F;
14'h1f9a:data=8'hFF;
14'h1f9b:data=8'hFF;
14'h1f9c:data=8'hFF;
14'h1f9d:data=8'hFF;
14'h1f9e:data=8'hFF;
14'h1f9f:data=8'hFF;
14'h1fa0:data=8'hFF;
14'h1fa1:data=8'hFF;
14'h1fa2:data=8'hFF;
14'h1fa3:data=8'hFF;
14'h1fa4:data=8'hFF;
14'h1fa5:data=8'hFC;
14'h1fa6:data=8'h00;
14'h1fa7:data=8'h00;
14'h1fc0:data=8'h00;
14'h1fc1:data=8'h03;
14'h1fc2:data=8'hFF;
14'h1fc3:data=8'hFE;
14'h1fc4:data=8'h00;
14'h1fc5:data=8'h00;
14'h1fc6:data=8'h00;
14'h1fc7:data=8'h00;
14'h1fc8:data=8'h00;
14'h1fc9:data=8'h1F;
14'h1fca:data=8'hFF;
14'h1fcb:data=8'hFF;
14'h1fcc:data=8'hF8;
14'h1fcd:data=8'h00;
14'h1fce:data=8'h00;
14'h1fcf:data=8'h00;
14'h1fd0:data=8'h00;
14'h1fd1:data=8'h07;
14'h1fd2:data=8'hFF;
14'h1fd3:data=8'hFF;
14'h1fd4:data=8'hFC;
14'h1fd5:data=8'h00;
14'h1fd6:data=8'h00;
14'h1fd7:data=8'h00;
14'h1fd8:data=8'h00;
14'h1fd9:data=8'h1F;
14'h1fda:data=8'hFF;
14'h1fdb:data=8'hFF;
14'h1fdc:data=8'hFF;
14'h1fdd:data=8'hFF;
14'h1fde:data=8'hFF;
14'h1fdf:data=8'hFF;
14'h1fe0:data=8'hFF;
14'h1fe1:data=8'hFF;
14'h1fe2:data=8'hFF;
14'h1fe3:data=8'hFF;
14'h1fe4:data=8'hFF;
14'h1fe5:data=8'hFC;
14'h1fe6:data=8'h00;
14'h1fe7:data=8'h00;
14'h2000:data=8'h00;
14'h2001:data=8'h03;
14'h2002:data=8'hFF;
14'h2003:data=8'hFE;
14'h2004:data=8'h00;
14'h2005:data=8'h00;
14'h2006:data=8'h00;
14'h2007:data=8'h00;
14'h2008:data=8'h00;
14'h2009:data=8'h1F;
14'h200a:data=8'hFF;
14'h200b:data=8'hFF;
14'h200c:data=8'hF8;
14'h200d:data=8'h00;
14'h200e:data=8'h00;
14'h200f:data=8'h00;
14'h2010:data=8'h00;
14'h2011:data=8'h07;
14'h2012:data=8'hFF;
14'h2013:data=8'hFF;
14'h2014:data=8'hFC;
14'h2015:data=8'h00;
14'h2016:data=8'h00;
14'h2017:data=8'h00;
14'h2018:data=8'h00;
14'h2019:data=8'h1F;
14'h201a:data=8'hFF;
14'h201b:data=8'hFF;
14'h201c:data=8'hFF;
14'h201d:data=8'hFF;
14'h201e:data=8'hFF;
14'h201f:data=8'hFF;
14'h2020:data=8'hFF;
14'h2021:data=8'hFF;
14'h2022:data=8'hFF;
14'h2023:data=8'hFF;
14'h2024:data=8'hFF;
14'h2025:data=8'hFC;
14'h2026:data=8'h00;
14'h2027:data=8'h00;
14'h2040:data=8'h00;
14'h2041:data=8'h03;
14'h2042:data=8'hFF;
14'h2043:data=8'hFE;
14'h2044:data=8'h00;
14'h2045:data=8'h00;
14'h2046:data=8'h00;
14'h2047:data=8'h00;
14'h2048:data=8'h00;
14'h2049:data=8'h1F;
14'h204a:data=8'hFF;
14'h204b:data=8'hFF;
14'h204c:data=8'hF8;
14'h204d:data=8'h00;
14'h204e:data=8'h00;
14'h204f:data=8'h00;
14'h2050:data=8'h00;
14'h2051:data=8'h07;
14'h2052:data=8'hFF;
14'h2053:data=8'hFF;
14'h2054:data=8'hFC;
14'h2055:data=8'h00;
14'h2056:data=8'h00;
14'h2057:data=8'h00;
14'h2058:data=8'h00;
14'h2059:data=8'h1F;
14'h205a:data=8'hFF;
14'h205b:data=8'hFF;
14'h205c:data=8'hFF;
14'h205d:data=8'hFF;
14'h205e:data=8'hFF;
14'h205f:data=8'hFF;
14'h2060:data=8'hFF;
14'h2061:data=8'hFF;
14'h2062:data=8'hFF;
14'h2063:data=8'hFF;
14'h2064:data=8'hFF;
14'h2065:data=8'hFC;
14'h2066:data=8'h00;
14'h2067:data=8'h00;
14'h2080:data=8'h00;
14'h2081:data=8'h03;
14'h2082:data=8'hFF;
14'h2083:data=8'hFE;
14'h2084:data=8'h00;
14'h2085:data=8'h00;
14'h2086:data=8'h00;
14'h2087:data=8'h00;
14'h2088:data=8'h00;
14'h2089:data=8'h1F;
14'h208a:data=8'hFF;
14'h208b:data=8'hFF;
14'h208c:data=8'hF8;
14'h208d:data=8'h00;
14'h208e:data=8'h00;
14'h208f:data=8'h00;
14'h2090:data=8'h00;
14'h2091:data=8'h07;
14'h2092:data=8'hFF;
14'h2093:data=8'hFF;
14'h2094:data=8'hFC;
14'h2095:data=8'h00;
14'h2096:data=8'h00;
14'h2097:data=8'h00;
14'h2098:data=8'h00;
14'h2099:data=8'h1F;
14'h209a:data=8'hFF;
14'h209b:data=8'hFF;
14'h209c:data=8'hFF;
14'h209d:data=8'hFF;
14'h209e:data=8'hFF;
14'h209f:data=8'hFF;
14'h20a0:data=8'hFF;
14'h20a1:data=8'hFF;
14'h20a2:data=8'hFF;
14'h20a3:data=8'hFF;
14'h20a4:data=8'hFF;
14'h20a5:data=8'hFC;
14'h20a6:data=8'h00;
14'h20a7:data=8'h00;
14'h20c0:data=8'h00;
14'h20c1:data=8'h03;
14'h20c2:data=8'hFF;
14'h20c3:data=8'hFF;
14'h20c4:data=8'h00;
14'h20c5:data=8'h00;
14'h20c6:data=8'h00;
14'h20c7:data=8'h00;
14'h20c8:data=8'h00;
14'h20c9:data=8'h1F;
14'h20ca:data=8'hFF;
14'h20cb:data=8'hFF;
14'h20cc:data=8'hF8;
14'h20cd:data=8'h00;
14'h20ce:data=8'h00;
14'h20cf:data=8'h00;
14'h20d0:data=8'h00;
14'h20d1:data=8'h07;
14'h20d2:data=8'hFF;
14'h20d3:data=8'hFF;
14'h20d4:data=8'hFC;
14'h20d5:data=8'h00;
14'h20d6:data=8'h00;
14'h20d7:data=8'h00;
14'h20d8:data=8'h00;
14'h20d9:data=8'h1F;
14'h20da:data=8'hFF;
14'h20db:data=8'hFF;
14'h20dc:data=8'hFF;
14'h20dd:data=8'hFF;
14'h20de:data=8'hFF;
14'h20df:data=8'hFF;
14'h20e0:data=8'hFF;
14'h20e1:data=8'hFF;
14'h20e2:data=8'hFF;
14'h20e3:data=8'hFF;
14'h20e4:data=8'hFF;
14'h20e5:data=8'hFC;
14'h20e6:data=8'h00;
14'h20e7:data=8'h00;
14'h2100:data=8'h00;
14'h2101:data=8'h03;
14'h2102:data=8'hFF;
14'h2103:data=8'hFF;
14'h2104:data=8'h00;
14'h2105:data=8'h00;
14'h2106:data=8'h00;
14'h2107:data=8'h00;
14'h2108:data=8'h00;
14'h2109:data=8'h1F;
14'h210a:data=8'hFF;
14'h210b:data=8'hFF;
14'h210c:data=8'hF8;
14'h210d:data=8'h00;
14'h210e:data=8'h00;
14'h210f:data=8'h00;
14'h2110:data=8'h00;
14'h2111:data=8'h07;
14'h2112:data=8'hFF;
14'h2113:data=8'hFF;
14'h2114:data=8'hFC;
14'h2115:data=8'h00;
14'h2116:data=8'h00;
14'h2117:data=8'h00;
14'h2118:data=8'h00;
14'h2119:data=8'h1F;
14'h211a:data=8'hFF;
14'h211b:data=8'hFF;
14'h211c:data=8'hFF;
14'h211d:data=8'hFF;
14'h211e:data=8'hFF;
14'h211f:data=8'hFF;
14'h2120:data=8'hFF;
14'h2121:data=8'hFF;
14'h2122:data=8'hFF;
14'h2123:data=8'hFF;
14'h2124:data=8'hFF;
14'h2125:data=8'hFC;
14'h2126:data=8'h00;
14'h2127:data=8'h00;
14'h2140:data=8'h00;
14'h2141:data=8'h03;
14'h2142:data=8'hFF;
14'h2143:data=8'hFF;
14'h2144:data=8'h00;
14'h2145:data=8'h00;
14'h2146:data=8'h00;
14'h2147:data=8'h00;
14'h2148:data=8'h00;
14'h2149:data=8'h1F;
14'h214a:data=8'hFF;
14'h214b:data=8'hFF;
14'h214c:data=8'hF8;
14'h214d:data=8'h00;
14'h214e:data=8'h00;
14'h214f:data=8'h00;
14'h2150:data=8'h00;
14'h2151:data=8'h07;
14'h2152:data=8'hFF;
14'h2153:data=8'hFF;
14'h2154:data=8'hFC;
14'h2155:data=8'h00;
14'h2156:data=8'h00;
14'h2157:data=8'h00;
14'h2158:data=8'h00;
14'h2159:data=8'h1F;
14'h215a:data=8'hFF;
14'h215b:data=8'hFF;
14'h215c:data=8'hFF;
14'h215d:data=8'hFF;
14'h215e:data=8'hFF;
14'h215f:data=8'hFF;
14'h2160:data=8'hFF;
14'h2161:data=8'hFF;
14'h2162:data=8'hFF;
14'h2163:data=8'hFF;
14'h2164:data=8'hFF;
14'h2165:data=8'hFC;
14'h2166:data=8'h00;
14'h2167:data=8'h00;
14'h2180:data=8'h00;
14'h2181:data=8'h03;
14'h2182:data=8'hFF;
14'h2183:data=8'hFF;
14'h2184:data=8'h00;
14'h2185:data=8'h00;
14'h2186:data=8'h00;
14'h2187:data=8'h00;
14'h2188:data=8'h00;
14'h2189:data=8'h1F;
14'h218a:data=8'hFF;
14'h218b:data=8'hFF;
14'h218c:data=8'hF8;
14'h218d:data=8'h00;
14'h218e:data=8'h00;
14'h218f:data=8'h00;
14'h2190:data=8'h00;
14'h2191:data=8'h07;
14'h2192:data=8'hFF;
14'h2193:data=8'hFF;
14'h2194:data=8'hFC;
14'h2195:data=8'h00;
14'h2196:data=8'h00;
14'h2197:data=8'h00;
14'h2198:data=8'h00;
14'h2199:data=8'h1F;
14'h219a:data=8'hFF;
14'h219b:data=8'hFF;
14'h219c:data=8'hFF;
14'h219d:data=8'hFF;
14'h219e:data=8'hFF;
14'h219f:data=8'hFF;
14'h21a0:data=8'hFF;
14'h21a1:data=8'hFF;
14'h21a2:data=8'hFF;
14'h21a3:data=8'hFF;
14'h21a4:data=8'hFF;
14'h21a5:data=8'hFC;
14'h21a6:data=8'h00;
14'h21a7:data=8'h00;
14'h21c0:data=8'h00;
14'h21c1:data=8'h03;
14'h21c2:data=8'hFF;
14'h21c3:data=8'hFF;
14'h21c4:data=8'h00;
14'h21c5:data=8'h00;
14'h21c6:data=8'h00;
14'h21c7:data=8'h00;
14'h21c8:data=8'h00;
14'h21c9:data=8'h1F;
14'h21ca:data=8'hFF;
14'h21cb:data=8'hFF;
14'h21cc:data=8'hF8;
14'h21cd:data=8'h00;
14'h21ce:data=8'h00;
14'h21cf:data=8'h00;
14'h21d0:data=8'h00;
14'h21d1:data=8'h07;
14'h21d2:data=8'hFF;
14'h21d3:data=8'hFF;
14'h21d4:data=8'hFC;
14'h21d5:data=8'h00;
14'h21d6:data=8'h00;
14'h21d7:data=8'h00;
14'h21d8:data=8'h00;
14'h21d9:data=8'h1F;
14'h21da:data=8'hFF;
14'h21db:data=8'hFF;
14'h21dc:data=8'hFF;
14'h21dd:data=8'hFF;
14'h21de:data=8'hFF;
14'h21df:data=8'hFF;
14'h21e0:data=8'hFF;
14'h21e1:data=8'hFF;
14'h21e2:data=8'hFF;
14'h21e3:data=8'hFF;
14'h21e4:data=8'hFF;
14'h21e5:data=8'hFC;
14'h21e6:data=8'h00;
14'h21e7:data=8'h00;
14'h2200:data=8'h00;
14'h2201:data=8'h03;
14'h2202:data=8'hFF;
14'h2203:data=8'hFF;
14'h2204:data=8'h00;
14'h2205:data=8'h00;
14'h2206:data=8'h00;
14'h2207:data=8'h00;
14'h2208:data=8'h00;
14'h2209:data=8'h1F;
14'h220a:data=8'hFF;
14'h220b:data=8'hFF;
14'h220c:data=8'hF8;
14'h220d:data=8'h00;
14'h220e:data=8'h00;
14'h220f:data=8'h00;
14'h2210:data=8'h00;
14'h2211:data=8'h07;
14'h2212:data=8'hFF;
14'h2213:data=8'hFF;
14'h2214:data=8'hFC;
14'h2215:data=8'h00;
14'h2216:data=8'h00;
14'h2217:data=8'h00;
14'h2218:data=8'h00;
14'h2219:data=8'h1F;
14'h221a:data=8'hFF;
14'h221b:data=8'hFF;
14'h221c:data=8'hFF;
14'h221d:data=8'hFF;
14'h221e:data=8'hFF;
14'h221f:data=8'hFF;
14'h2220:data=8'hFF;
14'h2221:data=8'hFF;
14'h2222:data=8'hFF;
14'h2223:data=8'hFF;
14'h2224:data=8'hFF;
14'h2225:data=8'hFC;
14'h2226:data=8'h00;
14'h2227:data=8'h00;
14'h2240:data=8'h00;
14'h2241:data=8'h03;
14'h2242:data=8'hFF;
14'h2243:data=8'hFF;
14'h2244:data=8'h00;
14'h2245:data=8'h00;
14'h2246:data=8'h00;
14'h2247:data=8'h00;
14'h2248:data=8'h00;
14'h2249:data=8'h1F;
14'h224a:data=8'hFF;
14'h224b:data=8'hFF;
14'h224c:data=8'hF8;
14'h224d:data=8'h00;
14'h224e:data=8'h00;
14'h224f:data=8'h00;
14'h2250:data=8'h00;
14'h2251:data=8'h07;
14'h2252:data=8'hFF;
14'h2253:data=8'hFF;
14'h2254:data=8'hFC;
14'h2255:data=8'h00;
14'h2256:data=8'h00;
14'h2257:data=8'h00;
14'h2258:data=8'h00;
14'h2259:data=8'h1F;
14'h225a:data=8'hFF;
14'h225b:data=8'hFF;
14'h225c:data=8'hFF;
14'h225d:data=8'hFF;
14'h225e:data=8'hFF;
14'h225f:data=8'hFF;
14'h2260:data=8'hFF;
14'h2261:data=8'hFF;
14'h2262:data=8'hFF;
14'h2263:data=8'hFF;
14'h2264:data=8'hFF;
14'h2265:data=8'hFC;
14'h2266:data=8'h00;
14'h2267:data=8'h00;
14'h2280:data=8'h00;
14'h2281:data=8'h03;
14'h2282:data=8'hFF;
14'h2283:data=8'hFF;
14'h2284:data=8'h00;
14'h2285:data=8'h00;
14'h2286:data=8'h00;
14'h2287:data=8'h00;
14'h2288:data=8'h00;
14'h2289:data=8'h1F;
14'h228a:data=8'hFF;
14'h228b:data=8'hFF;
14'h228c:data=8'hF8;
14'h228d:data=8'h00;
14'h228e:data=8'h00;
14'h228f:data=8'h00;
14'h2290:data=8'h00;
14'h2291:data=8'h07;
14'h2292:data=8'hFF;
14'h2293:data=8'hFF;
14'h2294:data=8'hFC;
14'h2295:data=8'h00;
14'h2296:data=8'h00;
14'h2297:data=8'h00;
14'h2298:data=8'h00;
14'h2299:data=8'h1F;
14'h229a:data=8'hFF;
14'h229b:data=8'hFF;
14'h229c:data=8'hFF;
14'h229d:data=8'hFF;
14'h229e:data=8'hFF;
14'h229f:data=8'hFF;
14'h22a0:data=8'hFF;
14'h22a1:data=8'hFF;
14'h22a2:data=8'hFF;
14'h22a3:data=8'hFF;
14'h22a4:data=8'hFF;
14'h22a5:data=8'hFC;
14'h22a6:data=8'h00;
14'h22a7:data=8'h00;
14'h22c0:data=8'h00;
14'h22c1:data=8'h03;
14'h22c2:data=8'hFF;
14'h22c3:data=8'hFF;
14'h22c4:data=8'h00;
14'h22c5:data=8'h00;
14'h22c6:data=8'h00;
14'h22c7:data=8'h00;
14'h22c8:data=8'h00;
14'h22c9:data=8'h1F;
14'h22ca:data=8'hFF;
14'h22cb:data=8'hFF;
14'h22cc:data=8'hF8;
14'h22cd:data=8'h00;
14'h22ce:data=8'h00;
14'h22cf:data=8'h00;
14'h22d0:data=8'h00;
14'h22d1:data=8'h07;
14'h22d2:data=8'hFF;
14'h22d3:data=8'hFF;
14'h22d4:data=8'hFC;
14'h22d5:data=8'h00;
14'h22d6:data=8'h00;
14'h22d7:data=8'h00;
14'h22d8:data=8'h00;
14'h22d9:data=8'h1F;
14'h22da:data=8'hFF;
14'h22db:data=8'hFF;
14'h22dc:data=8'hFF;
14'h22dd:data=8'hFF;
14'h22de:data=8'hFF;
14'h22df:data=8'hFF;
14'h22e0:data=8'hFF;
14'h22e1:data=8'hFF;
14'h22e2:data=8'hFF;
14'h22e3:data=8'hFF;
14'h22e4:data=8'hFF;
14'h22e5:data=8'hFC;
14'h22e6:data=8'h00;
14'h22e7:data=8'h00;
14'h2300:data=8'h00;
14'h2301:data=8'h03;
14'h2302:data=8'hFF;
14'h2303:data=8'hFF;
14'h2304:data=8'h00;
14'h2305:data=8'h00;
14'h2306:data=8'h00;
14'h2307:data=8'h00;
14'h2308:data=8'h00;
14'h2309:data=8'h1F;
14'h230a:data=8'hFF;
14'h230b:data=8'hFF;
14'h230c:data=8'hF8;
14'h230d:data=8'h00;
14'h230e:data=8'h00;
14'h230f:data=8'h00;
14'h2310:data=8'h00;
14'h2311:data=8'h07;
14'h2312:data=8'hFF;
14'h2313:data=8'hFF;
14'h2314:data=8'hFC;
14'h2315:data=8'h00;
14'h2316:data=8'h00;
14'h2317:data=8'h00;
14'h2318:data=8'h00;
14'h2319:data=8'h00;
14'h231a:data=8'h3F;
14'h231b:data=8'hFF;
14'h231c:data=8'hFF;
14'h231d:data=8'hFF;
14'h231e:data=8'hFF;
14'h231f:data=8'hFF;
14'h2320:data=8'hFF;
14'h2321:data=8'hFF;
14'h2322:data=8'hC0;
14'h2323:data=8'h00;
14'h2324:data=8'h00;
14'h2325:data=8'h00;
14'h2326:data=8'h00;
14'h2327:data=8'h00;
14'h2340:data=8'h00;
14'h2341:data=8'h03;
14'h2342:data=8'hFF;
14'h2343:data=8'hFF;
14'h2344:data=8'h00;
14'h2345:data=8'h00;
14'h2346:data=8'h00;
14'h2347:data=8'h00;
14'h2348:data=8'h00;
14'h2349:data=8'h1F;
14'h234a:data=8'hFF;
14'h234b:data=8'hFF;
14'h234c:data=8'hF8;
14'h234d:data=8'h00;
14'h234e:data=8'h00;
14'h234f:data=8'h00;
14'h2350:data=8'h00;
14'h2351:data=8'h07;
14'h2352:data=8'hFF;
14'h2353:data=8'hFF;
14'h2354:data=8'hFC;
14'h2355:data=8'h00;
14'h2356:data=8'h00;
14'h2357:data=8'h00;
14'h2358:data=8'h00;
14'h2359:data=8'h00;
14'h235a:data=8'h3F;
14'h235b:data=8'hFF;
14'h235c:data=8'hFF;
14'h235d:data=8'hFF;
14'h235e:data=8'hFF;
14'h235f:data=8'hFF;
14'h2360:data=8'hFF;
14'h2361:data=8'hFE;
14'h2362:data=8'h00;
14'h2363:data=8'h00;
14'h2364:data=8'h00;
14'h2365:data=8'h00;
14'h2366:data=8'h00;
14'h2367:data=8'h00;
14'h2380:data=8'h00;
14'h2381:data=8'h03;
14'h2382:data=8'hFF;
14'h2383:data=8'hFF;
14'h2384:data=8'h00;
14'h2385:data=8'h00;
14'h2386:data=8'h00;
14'h2387:data=8'h00;
14'h2388:data=8'h00;
14'h2389:data=8'h1F;
14'h238a:data=8'hFF;
14'h238b:data=8'hFF;
14'h238c:data=8'hF8;
14'h238d:data=8'h00;
14'h238e:data=8'h00;
14'h238f:data=8'h00;
14'h2390:data=8'h00;
14'h2391:data=8'h07;
14'h2392:data=8'hFF;
14'h2393:data=8'hFF;
14'h2394:data=8'hFC;
14'h2395:data=8'h00;
14'h2396:data=8'h00;
14'h2397:data=8'h00;
14'h2398:data=8'h00;
14'h2399:data=8'h00;
14'h239a:data=8'h3F;
14'h239b:data=8'hFF;
14'h239c:data=8'hFF;
14'h239d:data=8'hFF;
14'h239e:data=8'hFF;
14'h239f:data=8'hFF;
14'h23a0:data=8'hFF;
14'h23a1:data=8'hF0;
14'h23a2:data=8'h00;
14'h23a3:data=8'h00;
14'h23a4:data=8'h00;
14'h23a5:data=8'h00;
14'h23a6:data=8'h00;
14'h23a7:data=8'h00;
14'h23c0:data=8'h00;
14'h23c1:data=8'h03;
14'h23c2:data=8'hFF;
14'h23c3:data=8'hFF;
14'h23c4:data=8'h00;
14'h23c5:data=8'h00;
14'h23c6:data=8'h00;
14'h23c7:data=8'h00;
14'h23c8:data=8'h00;
14'h23c9:data=8'h1F;
14'h23ca:data=8'hFF;
14'h23cb:data=8'hFF;
14'h23cc:data=8'hF8;
14'h23cd:data=8'h00;
14'h23ce:data=8'h00;
14'h23cf:data=8'h00;
14'h23d0:data=8'h00;
14'h23d1:data=8'h07;
14'h23d2:data=8'hFF;
14'h23d3:data=8'hFF;
14'h23d4:data=8'hFE;
14'h23d5:data=8'h00;
14'h23d6:data=8'h00;
14'h23d7:data=8'h00;
14'h23d8:data=8'h00;
14'h23d9:data=8'h00;
14'h23da:data=8'h3F;
14'h23db:data=8'hFF;
14'h23dc:data=8'hFF;
14'h23dd:data=8'hFF;
14'h23de:data=8'hFF;
14'h23df:data=8'hFF;
14'h23e0:data=8'hFF;
14'h23e1:data=8'h80;
14'h23e2:data=8'h00;
14'h23e3:data=8'h00;
14'h23e4:data=8'h00;
14'h23e5:data=8'h00;
14'h23e6:data=8'h00;
14'h23e7:data=8'h00;
14'h2400:data=8'h00;
14'h2401:data=8'h03;
14'h2402:data=8'hFF;
14'h2403:data=8'hFF;
14'h2404:data=8'h00;
14'h2405:data=8'h00;
14'h2406:data=8'h00;
14'h2407:data=8'h00;
14'h2408:data=8'h00;
14'h2409:data=8'h1F;
14'h240a:data=8'hFF;
14'h240b:data=8'hFF;
14'h240c:data=8'hF8;
14'h240d:data=8'h00;
14'h240e:data=8'h00;
14'h240f:data=8'h00;
14'h2410:data=8'h00;
14'h2411:data=8'h07;
14'h2412:data=8'hFF;
14'h2413:data=8'hFF;
14'h2414:data=8'hFE;
14'h2415:data=8'h00;
14'h2416:data=8'h00;
14'h2417:data=8'h00;
14'h2418:data=8'h00;
14'h2419:data=8'h00;
14'h241a:data=8'h3F;
14'h241b:data=8'hFF;
14'h241c:data=8'hFF;
14'h241d:data=8'hFF;
14'h241e:data=8'hFF;
14'h241f:data=8'hFF;
14'h2420:data=8'hFC;
14'h2421:data=8'h00;
14'h2422:data=8'h00;
14'h2423:data=8'h00;
14'h2424:data=8'h00;
14'h2425:data=8'h00;
14'h2426:data=8'h00;
14'h2427:data=8'h00;
14'h2440:data=8'h00;
14'h2441:data=8'h03;
14'h2442:data=8'hFF;
14'h2443:data=8'hFF;
14'h2444:data=8'h00;
14'h2445:data=8'h00;
14'h2446:data=8'h00;
14'h2447:data=8'h00;
14'h2448:data=8'h00;
14'h2449:data=8'h1F;
14'h244a:data=8'hFF;
14'h244b:data=8'hFF;
14'h244c:data=8'hF8;
14'h244d:data=8'h00;
14'h244e:data=8'h00;
14'h244f:data=8'h00;
14'h2450:data=8'h00;
14'h2451:data=8'h07;
14'h2452:data=8'hFF;
14'h2453:data=8'hFF;
14'h2454:data=8'hFE;
14'h2455:data=8'h00;
14'h2456:data=8'h00;
14'h2457:data=8'h00;
14'h2458:data=8'h00;
14'h2459:data=8'h00;
14'h245a:data=8'h3F;
14'h245b:data=8'hFF;
14'h245c:data=8'hFF;
14'h245d:data=8'hFF;
14'h245e:data=8'hFF;
14'h245f:data=8'hFF;
14'h2460:data=8'hC0;
14'h2461:data=8'h00;
14'h2462:data=8'h00;
14'h2463:data=8'h00;
14'h2464:data=8'h00;
14'h2465:data=8'h00;
14'h2466:data=8'h00;
14'h2467:data=8'h03;
14'h2480:data=8'h00;
14'h2481:data=8'h01;
14'h2482:data=8'hFF;
14'h2483:data=8'hFF;
14'h2484:data=8'h00;
14'h2485:data=8'h00;
14'h2486:data=8'h00;
14'h2487:data=8'h00;
14'h2488:data=8'h00;
14'h2489:data=8'h1F;
14'h248a:data=8'hFF;
14'h248b:data=8'hFF;
14'h248c:data=8'hF8;
14'h248d:data=8'h00;
14'h248e:data=8'h00;
14'h248f:data=8'h00;
14'h2490:data=8'h00;
14'h2491:data=8'h07;
14'h2492:data=8'hFF;
14'h2493:data=8'hFF;
14'h2494:data=8'hFE;
14'h2495:data=8'h00;
14'h2496:data=8'h00;
14'h2497:data=8'h00;
14'h2498:data=8'h00;
14'h2499:data=8'h00;
14'h249a:data=8'h3F;
14'h249b:data=8'hFF;
14'h249c:data=8'hFF;
14'h249d:data=8'hFF;
14'h249e:data=8'hFF;
14'h249f:data=8'hFE;
14'h24a0:data=8'h00;
14'h24a1:data=8'h00;
14'h24a2:data=8'h00;
14'h24a3:data=8'h00;
14'h24a4:data=8'h00;
14'h24a5:data=8'h00;
14'h24a6:data=8'h00;
14'h24a7:data=8'h1C;
14'h24c0:data=8'h00;
14'h24c1:data=8'h01;
14'h24c2:data=8'hFF;
14'h24c3:data=8'hFF;
14'h24c4:data=8'h00;
14'h24c5:data=8'h00;
14'h24c6:data=8'h00;
14'h24c7:data=8'h00;
14'h24c8:data=8'h00;
14'h24c9:data=8'h1F;
14'h24ca:data=8'hFF;
14'h24cb:data=8'hFF;
14'h24cc:data=8'hF8;
14'h24cd:data=8'h00;
14'h24ce:data=8'h00;
14'h24cf:data=8'h00;
14'h24d0:data=8'h00;
14'h24d1:data=8'h07;
14'h24d2:data=8'hFF;
14'h24d3:data=8'hFF;
14'h24d4:data=8'hFE;
14'h24d5:data=8'h00;
14'h24d6:data=8'h00;
14'h24d7:data=8'h00;
14'h24d8:data=8'h00;
14'h24d9:data=8'h00;
14'h24da:data=8'h3F;
14'h24db:data=8'hFF;
14'h24dc:data=8'hFF;
14'h24dd:data=8'hFF;
14'h24de:data=8'hFF;
14'h24df:data=8'hF0;
14'h24e0:data=8'h00;
14'h24e1:data=8'h00;
14'h24e2:data=8'h00;
14'h24e3:data=8'h00;
14'h24e4:data=8'h00;
14'h24e5:data=8'h00;
14'h24e6:data=8'h00;
14'h24e7:data=8'hE0;
14'h2500:data=8'h00;
14'h2501:data=8'h01;
14'h2502:data=8'hFF;
14'h2503:data=8'hFF;
14'h2504:data=8'h00;
14'h2505:data=8'h00;
14'h2506:data=8'h00;
14'h2507:data=8'h00;
14'h2508:data=8'h00;
14'h2509:data=8'h1F;
14'h250a:data=8'hFF;
14'h250b:data=8'hFF;
14'h250c:data=8'hF8;
14'h250d:data=8'h00;
14'h250e:data=8'h00;
14'h250f:data=8'h00;
14'h2510:data=8'h00;
14'h2511:data=8'h07;
14'h2512:data=8'hFF;
14'h2513:data=8'hFF;
14'h2514:data=8'hFE;
14'h2515:data=8'h00;
14'h2516:data=8'h00;
14'h2517:data=8'h00;
14'h2518:data=8'h00;
14'h2519:data=8'h00;
14'h251a:data=8'h3F;
14'h251b:data=8'hFF;
14'h251c:data=8'hFF;
14'h251d:data=8'hFF;
14'h251e:data=8'hFF;
14'h251f:data=8'h80;
14'h2520:data=8'h00;
14'h2521:data=8'h00;
14'h2522:data=8'h00;
14'h2523:data=8'h00;
14'h2524:data=8'h00;
14'h2525:data=8'h00;
14'h2526:data=8'h07;
14'h2527:data=8'h00;
14'h2540:data=8'h00;
14'h2541:data=8'h01;
14'h2542:data=8'hFF;
14'h2543:data=8'hFF;
14'h2544:data=8'h00;
14'h2545:data=8'h00;
14'h2546:data=8'h00;
14'h2547:data=8'h00;
14'h2548:data=8'h00;
14'h2549:data=8'h1F;
14'h254a:data=8'hFF;
14'h254b:data=8'hFF;
14'h254c:data=8'hF8;
14'h254d:data=8'h00;
14'h254e:data=8'h00;
14'h254f:data=8'h00;
14'h2550:data=8'h00;
14'h2551:data=8'h07;
14'h2552:data=8'hFF;
14'h2553:data=8'hFF;
14'h2554:data=8'hFE;
14'h2555:data=8'h00;
14'h2556:data=8'h00;
14'h2557:data=8'h00;
14'h2558:data=8'h00;
14'h2559:data=8'h00;
14'h255a:data=8'h3F;
14'h255b:data=8'hFF;
14'h255c:data=8'hFF;
14'h255d:data=8'hFF;
14'h255e:data=8'hFC;
14'h255f:data=8'h00;
14'h2560:data=8'h00;
14'h2561:data=8'h00;
14'h2562:data=8'h00;
14'h2563:data=8'h00;
14'h2564:data=8'h00;
14'h2565:data=8'h00;
14'h2566:data=8'h38;
14'h2567:data=8'h00;
14'h2580:data=8'h00;
14'h2581:data=8'h01;
14'h2582:data=8'hFF;
14'h2583:data=8'hFF;
14'h2584:data=8'h00;
14'h2585:data=8'h00;
14'h2586:data=8'h00;
14'h2587:data=8'h00;
14'h2588:data=8'h00;
14'h2589:data=8'h1F;
14'h258a:data=8'hFF;
14'h258b:data=8'hFF;
14'h258c:data=8'hF8;
14'h258d:data=8'h00;
14'h258e:data=8'h00;
14'h258f:data=8'h00;
14'h2590:data=8'h00;
14'h2591:data=8'h07;
14'h2592:data=8'hFF;
14'h2593:data=8'hFF;
14'h2594:data=8'hFE;
14'h2595:data=8'h00;
14'h2596:data=8'h00;
14'h2597:data=8'h00;
14'h2598:data=8'h00;
14'h2599:data=8'h00;
14'h259a:data=8'h3F;
14'h259b:data=8'hFF;
14'h259c:data=8'hFF;
14'h259d:data=8'hFF;
14'h259e:data=8'hE0;
14'h259f:data=8'h00;
14'h25a0:data=8'h00;
14'h25a1:data=8'h00;
14'h25a2:data=8'h00;
14'h25a3:data=8'h00;
14'h25a4:data=8'h00;
14'h25a5:data=8'h01;
14'h25a6:data=8'hC0;
14'h25a7:data=8'h00;
14'h25c0:data=8'h00;
14'h25c1:data=8'h01;
14'h25c2:data=8'hFF;
14'h25c3:data=8'hFF;
14'h25c4:data=8'h00;
14'h25c5:data=8'h00;
14'h25c6:data=8'h00;
14'h25c7:data=8'h00;
14'h25c8:data=8'h00;
14'h25c9:data=8'h1F;
14'h25ca:data=8'hFF;
14'h25cb:data=8'hFF;
14'h25cc:data=8'hF8;
14'h25cd:data=8'h00;
14'h25ce:data=8'h00;
14'h25cf:data=8'h00;
14'h25d0:data=8'h00;
14'h25d1:data=8'h07;
14'h25d2:data=8'hFF;
14'h25d3:data=8'hFF;
14'h25d4:data=8'hFE;
14'h25d5:data=8'h00;
14'h25d6:data=8'h00;
14'h25d7:data=8'h00;
14'h25d8:data=8'h00;
14'h25d9:data=8'h00;
14'h25da:data=8'h3F;
14'h25db:data=8'hFF;
14'h25dc:data=8'hFF;
14'h25dd:data=8'hFE;
14'h25de:data=8'h00;
14'h25df:data=8'h00;
14'h25e0:data=8'h00;
14'h25e1:data=8'h00;
14'h25e2:data=8'h00;
14'h25e3:data=8'h00;
14'h25e4:data=8'h00;
14'h25e5:data=8'h0E;
14'h25e6:data=8'h00;
14'h25e7:data=8'h00;
14'h2600:data=8'h00;
14'h2601:data=8'h01;
14'h2602:data=8'hFF;
14'h2603:data=8'hFF;
14'h2604:data=8'h00;
14'h2605:data=8'h00;
14'h2606:data=8'h00;
14'h2607:data=8'h00;
14'h2608:data=8'h00;
14'h2609:data=8'h1F;
14'h260a:data=8'hFF;
14'h260b:data=8'hFF;
14'h260c:data=8'hF8;
14'h260d:data=8'h00;
14'h260e:data=8'h00;
14'h260f:data=8'h00;
14'h2610:data=8'h00;
14'h2611:data=8'h07;
14'h2612:data=8'hFF;
14'h2613:data=8'hFF;
14'h2614:data=8'hFE;
14'h2615:data=8'h00;
14'h2616:data=8'h00;
14'h2617:data=8'h00;
14'h2618:data=8'h00;
14'h2619:data=8'h00;
14'h261a:data=8'h3F;
14'h261b:data=8'hFF;
14'h261c:data=8'hFF;
14'h261d:data=8'hF0;
14'h261e:data=8'h00;
14'h261f:data=8'h00;
14'h2620:data=8'h00;
14'h2621:data=8'h00;
14'h2622:data=8'h00;
14'h2623:data=8'h00;
14'h2624:data=8'h00;
14'h2625:data=8'h70;
14'h2626:data=8'h00;
14'h2627:data=8'h00;
14'h2640:data=8'h00;
14'h2641:data=8'h01;
14'h2642:data=8'hFF;
14'h2643:data=8'hFF;
14'h2644:data=8'h00;
14'h2645:data=8'h00;
14'h2646:data=8'h00;
14'h2647:data=8'h00;
14'h2648:data=8'h00;
14'h2649:data=8'h1F;
14'h264a:data=8'hFF;
14'h264b:data=8'hFF;
14'h264c:data=8'hF8;
14'h264d:data=8'h00;
14'h264e:data=8'h00;
14'h264f:data=8'h00;
14'h2650:data=8'h00;
14'h2651:data=8'h07;
14'h2652:data=8'hFF;
14'h2653:data=8'hFF;
14'h2654:data=8'hFE;
14'h2655:data=8'h00;
14'h2656:data=8'h00;
14'h2657:data=8'h00;
14'h2658:data=8'h00;
14'h2659:data=8'h00;
14'h265a:data=8'h3F;
14'h265b:data=8'hFF;
14'h265c:data=8'hFF;
14'h265d:data=8'h80;
14'h265e:data=8'h00;
14'h265f:data=8'h00;
14'h2660:data=8'h00;
14'h2661:data=8'h00;
14'h2662:data=8'h00;
14'h2663:data=8'h00;
14'h2664:data=8'h03;
14'h2665:data=8'h80;
14'h2666:data=8'h00;
14'h2667:data=8'h00;
14'h2680:data=8'h00;
14'h2681:data=8'h01;
14'h2682:data=8'hFF;
14'h2683:data=8'hFF;
14'h2684:data=8'h80;
14'h2685:data=8'h00;
14'h2686:data=8'h00;
14'h2687:data=8'h00;
14'h2688:data=8'h00;
14'h2689:data=8'h1F;
14'h268a:data=8'hFF;
14'h268b:data=8'hFF;
14'h268c:data=8'hF8;
14'h268d:data=8'h00;
14'h268e:data=8'h00;
14'h268f:data=8'h00;
14'h2690:data=8'h00;
14'h2691:data=8'h07;
14'h2692:data=8'hFF;
14'h2693:data=8'hFF;
14'h2694:data=8'hFE;
14'h2695:data=8'h00;
14'h2696:data=8'h00;
14'h2697:data=8'h00;
14'h2698:data=8'h00;
14'h2699:data=8'h00;
14'h269a:data=8'h3F;
14'h269b:data=8'hFF;
14'h269c:data=8'hFC;
14'h269d:data=8'h00;
14'h269e:data=8'h00;
14'h269f:data=8'h00;
14'h26a0:data=8'h00;
14'h26a1:data=8'h00;
14'h26a2:data=8'h00;
14'h26a3:data=8'h00;
14'h26a4:data=8'h1C;
14'h26a5:data=8'h00;
14'h26a6:data=8'h00;
14'h26a7:data=8'h00;
14'h26c0:data=8'h00;
14'h26c1:data=8'h01;
14'h26c2:data=8'hFF;
14'h26c3:data=8'hFF;
14'h26c4:data=8'h80;
14'h26c5:data=8'h00;
14'h26c6:data=8'h00;
14'h26c7:data=8'h00;
14'h26c8:data=8'h00;
14'h26c9:data=8'h1F;
14'h26ca:data=8'hFF;
14'h26cb:data=8'hFF;
14'h26cc:data=8'hF8;
14'h26cd:data=8'h00;
14'h26ce:data=8'h00;
14'h26cf:data=8'h00;
14'h26d0:data=8'h00;
14'h26d1:data=8'h07;
14'h26d2:data=8'hFF;
14'h26d3:data=8'hFF;
14'h26d4:data=8'hFE;
14'h26d5:data=8'h00;
14'h26d6:data=8'h00;
14'h26d7:data=8'h00;
14'h26d8:data=8'h00;
14'h26d9:data=8'h00;
14'h26da:data=8'h3F;
14'h26db:data=8'hFF;
14'h26dc:data=8'hC0;
14'h26dd:data=8'h00;
14'h26de:data=8'h00;
14'h26df:data=8'h00;
14'h26e0:data=8'h00;
14'h26e1:data=8'h00;
14'h26e2:data=8'h00;
14'h26e3:data=8'h00;
14'h26e4:data=8'hC0;
14'h26e5:data=8'h00;
14'h26e6:data=8'h00;
14'h26e7:data=8'h00;
14'h2700:data=8'h00;
14'h2701:data=8'h01;
14'h2702:data=8'hFF;
14'h2703:data=8'hFF;
14'h2704:data=8'h80;
14'h2705:data=8'h00;
14'h2706:data=8'h00;
14'h2707:data=8'h00;
14'h2708:data=8'h00;
14'h2709:data=8'h1F;
14'h270a:data=8'hFF;
14'h270b:data=8'hFF;
14'h270c:data=8'hF8;
14'h270d:data=8'h00;
14'h270e:data=8'h00;
14'h270f:data=8'h00;
14'h2710:data=8'h00;
14'h2711:data=8'h07;
14'h2712:data=8'hFF;
14'h2713:data=8'hFF;
14'h2714:data=8'hFE;
14'h2715:data=8'h00;
14'h2716:data=8'h00;
14'h2717:data=8'h00;
14'h2718:data=8'h00;
14'h2719:data=8'h00;
14'h271a:data=8'h3F;
14'h271b:data=8'hFE;
14'h271c:data=8'h00;
14'h271d:data=8'h00;
14'h271e:data=8'h00;
14'h271f:data=8'h00;
14'h2720:data=8'h00;
14'h2721:data=8'h00;
14'h2722:data=8'h00;
14'h2723:data=8'h06;
14'h2724:data=8'h00;
14'h2725:data=8'h00;
14'h2726:data=8'h00;
14'h2727:data=8'h00;
14'h2740:data=8'h00;
14'h2741:data=8'h01;
14'h2742:data=8'hFF;
14'h2743:data=8'hFF;
14'h2744:data=8'h80;
14'h2745:data=8'h00;
14'h2746:data=8'h00;
14'h2747:data=8'h00;
14'h2748:data=8'h00;
14'h2749:data=8'h1F;
14'h274a:data=8'hFF;
14'h274b:data=8'hFF;
14'h274c:data=8'hF8;
14'h274d:data=8'h00;
14'h274e:data=8'h00;
14'h274f:data=8'h00;
14'h2750:data=8'h00;
14'h2751:data=8'h07;
14'h2752:data=8'hFF;
14'h2753:data=8'hFF;
14'h2754:data=8'hFE;
14'h2755:data=8'h00;
14'h2756:data=8'h00;
14'h2757:data=8'h00;
14'h2758:data=8'h00;
14'h2759:data=8'h00;
14'h275a:data=8'h1F;
14'h275b:data=8'hF0;
14'h275c:data=8'h00;
14'h275d:data=8'h00;
14'h275e:data=8'h00;
14'h275f:data=8'h00;
14'h2760:data=8'h00;
14'h2761:data=8'h00;
14'h2762:data=8'h00;
14'h2763:data=8'h30;
14'h2764:data=8'h00;
14'h2765:data=8'h00;
14'h2766:data=8'h00;
14'h2767:data=8'h00;
14'h2780:data=8'h00;
14'h2781:data=8'h01;
14'h2782:data=8'hFF;
14'h2783:data=8'hFF;
14'h2784:data=8'h80;
14'h2785:data=8'h00;
14'h2786:data=8'h00;
14'h2787:data=8'h00;
14'h2788:data=8'h00;
14'h2789:data=8'h0F;
14'h278a:data=8'hFF;
14'h278b:data=8'hFF;
14'h278c:data=8'hF8;
14'h278d:data=8'h00;
14'h278e:data=8'h00;
14'h278f:data=8'h00;
14'h2790:data=8'h00;
14'h2791:data=8'h07;
14'h2792:data=8'hFF;
14'h2793:data=8'hFF;
14'h2794:data=8'hFE;
14'h2795:data=8'h00;
14'h2796:data=8'h00;
14'h2797:data=8'h00;
14'h2798:data=8'h00;
14'h2799:data=8'h00;
14'h279a:data=8'h1F;
14'h279b:data=8'h80;
14'h279c:data=8'h00;
14'h279d:data=8'h00;
14'h279e:data=8'h00;
14'h279f:data=8'h00;
14'h27a0:data=8'h00;
14'h27a1:data=8'h00;
14'h27a2:data=8'h01;
14'h27a3:data=8'h80;
14'h27a4:data=8'h00;
14'h27a5:data=8'h00;
14'h27a6:data=8'h00;
14'h27a7:data=8'h00;
14'h27c0:data=8'h00;
14'h27c1:data=8'h01;
14'h27c2:data=8'hFF;
14'h27c3:data=8'hFF;
14'h27c4:data=8'h80;
14'h27c5:data=8'h00;
14'h27c6:data=8'h00;
14'h27c7:data=8'h00;
14'h27c8:data=8'h00;
14'h27c9:data=8'h0F;
14'h27ca:data=8'hFF;
14'h27cb:data=8'hFF;
14'h27cc:data=8'hF8;
14'h27cd:data=8'h00;
14'h27ce:data=8'h00;
14'h27cf:data=8'h00;
14'h27d0:data=8'h00;
14'h27d1:data=8'h07;
14'h27d2:data=8'hFF;
14'h27d3:data=8'hFF;
14'h27d4:data=8'hFE;
14'h27d5:data=8'h00;
14'h27d6:data=8'h00;
14'h27d7:data=8'h00;
14'h27d8:data=8'h00;
14'h27d9:data=8'h00;
14'h27da:data=8'h00;
14'h27db:data=8'h00;
14'h27dc:data=8'h00;
14'h27dd:data=8'h00;
14'h27de:data=8'h00;
14'h27df:data=8'h00;
14'h27e0:data=8'h00;
14'h27e1:data=8'h00;
14'h27e2:data=8'h1C;
14'h27e3:data=8'h00;
14'h27e4:data=8'h00;
14'h27e5:data=8'h00;
14'h27e6:data=8'h00;
14'h27e7:data=8'h00;
14'h2800:data=8'h00;
14'h2801:data=8'h01;
14'h2802:data=8'hFF;
14'h2803:data=8'hFF;
14'h2804:data=8'h80;
14'h2805:data=8'h00;
14'h2806:data=8'h00;
14'h2807:data=8'h00;
14'h2808:data=8'h00;
14'h2809:data=8'h00;
14'h280a:data=8'h03;
14'h280b:data=8'hFF;
14'h280c:data=8'hF8;
14'h280d:data=8'h00;
14'h280e:data=8'h00;
14'h280f:data=8'h00;
14'h2810:data=8'h00;
14'h2811:data=8'h07;
14'h2812:data=8'hFF;
14'h2813:data=8'hFF;
14'h2814:data=8'hFE;
14'h2815:data=8'h00;
14'h2816:data=8'h00;
14'h2817:data=8'h00;
14'h2818:data=8'h00;
14'h2819:data=8'h00;
14'h281a:data=8'h00;
14'h281b:data=8'h00;
14'h281c:data=8'h00;
14'h281d:data=8'h00;
14'h281e:data=8'h00;
14'h281f:data=8'h00;
14'h2820:data=8'h00;
14'h2821:data=8'h00;
14'h2822:data=8'hE0;
14'h2823:data=8'h00;
14'h2824:data=8'h00;
14'h2825:data=8'h00;
14'h2826:data=8'h00;
14'h2827:data=8'h01;
14'h2840:data=8'h00;
14'h2841:data=8'h01;
14'h2842:data=8'hFF;
14'h2843:data=8'hFF;
14'h2844:data=8'h80;
14'h2845:data=8'h00;
14'h2846:data=8'h00;
14'h2847:data=8'h00;
14'h2848:data=8'h00;
14'h2849:data=8'h00;
14'h284a:data=8'h03;
14'h284b:data=8'hFF;
14'h284c:data=8'hF8;
14'h284d:data=8'h00;
14'h284e:data=8'h00;
14'h284f:data=8'h00;
14'h2850:data=8'h00;
14'h2851:data=8'h07;
14'h2852:data=8'hFF;
14'h2853:data=8'hFF;
14'h2854:data=8'hFE;
14'h2855:data=8'h00;
14'h2856:data=8'h00;
14'h2857:data=8'h00;
14'h2858:data=8'h00;
14'h2859:data=8'h00;
14'h285a:data=8'h00;
14'h285b:data=8'h00;
14'h285c:data=8'h00;
14'h285d:data=8'h00;
14'h285e:data=8'h00;
14'h285f:data=8'h00;
14'h2860:data=8'h00;
14'h2861:data=8'h07;
14'h2862:data=8'h00;
14'h2863:data=8'h00;
14'h2864:data=8'h00;
14'h2865:data=8'h00;
14'h2866:data=8'h00;
14'h2867:data=8'h0C;
14'h2880:data=8'h00;
14'h2881:data=8'h01;
14'h2882:data=8'hFF;
14'h2883:data=8'hFF;
14'h2884:data=8'h80;
14'h2885:data=8'h00;
14'h2886:data=8'h00;
14'h2887:data=8'h00;
14'h2888:data=8'h00;
14'h2889:data=8'h00;
14'h288a:data=8'h03;
14'h288b:data=8'hFF;
14'h288c:data=8'hF8;
14'h288d:data=8'h00;
14'h288e:data=8'h00;
14'h288f:data=8'h00;
14'h2890:data=8'h00;
14'h2891:data=8'h07;
14'h2892:data=8'hFF;
14'h2893:data=8'hFF;
14'h2894:data=8'h00;
14'h2895:data=8'h00;
14'h2896:data=8'h00;
14'h2897:data=8'h00;
14'h2898:data=8'h00;
14'h2899:data=8'h00;
14'h289a:data=8'h00;
14'h289b:data=8'h00;
14'h289c:data=8'h00;
14'h289d:data=8'h00;
14'h289e:data=8'h00;
14'h289f:data=8'h00;
14'h28a0:data=8'h00;
14'h28a1:data=8'h38;
14'h28a2:data=8'h00;
14'h28a3:data=8'h00;
14'h28a4:data=8'h00;
14'h28a5:data=8'h00;
14'h28a6:data=8'h00;
14'h28a7:data=8'h60;
14'h28c0:data=8'h00;
14'h28c1:data=8'h01;
14'h28c2:data=8'hFF;
14'h28c3:data=8'hFF;
14'h28c4:data=8'h80;
14'h28c5:data=8'h00;
14'h28c6:data=8'h00;
14'h28c7:data=8'h00;
14'h28c8:data=8'h00;
14'h28c9:data=8'h00;
14'h28ca:data=8'h03;
14'h28cb:data=8'hFF;
14'h28cc:data=8'hFF;
14'h28cd:data=8'hFF;
14'h28ce:data=8'hFF;
14'h28cf:data=8'hFF;
14'h28d0:data=8'hFF;
14'h28d1:data=8'hFF;
14'h28d2:data=8'hFF;
14'h28d3:data=8'hFF;
14'h28d4:data=8'h00;
14'h28d5:data=8'h00;
14'h28d6:data=8'h00;
14'h28d7:data=8'h00;
14'h28d8:data=8'h00;
14'h28d9:data=8'h00;
14'h28da:data=8'h00;
14'h28db:data=8'h00;
14'h28dc:data=8'h00;
14'h28dd:data=8'h00;
14'h28de:data=8'h00;
14'h28df:data=8'h00;
14'h28e0:data=8'h01;
14'h28e1:data=8'hC0;
14'h28e2:data=8'h00;
14'h28e3:data=8'h00;
14'h28e4:data=8'h00;
14'h28e5:data=8'h00;
14'h28e6:data=8'h07;
14'h28e7:data=8'h00;
14'h2900:data=8'h00;
14'h2901:data=8'h01;
14'h2902:data=8'hFF;
14'h2903:data=8'hFF;
14'h2904:data=8'h80;
14'h2905:data=8'h00;
14'h2906:data=8'h00;
14'h2907:data=8'h00;
14'h2908:data=8'h00;
14'h2909:data=8'h00;
14'h290a:data=8'h03;
14'h290b:data=8'hFF;
14'h290c:data=8'hFF;
14'h290d:data=8'hFF;
14'h290e:data=8'hFF;
14'h290f:data=8'hFF;
14'h2910:data=8'hFF;
14'h2911:data=8'hFF;
14'h2912:data=8'hFF;
14'h2913:data=8'hFF;
14'h2914:data=8'h00;
14'h2915:data=8'h00;
14'h2916:data=8'h00;
14'h2917:data=8'h00;
14'h2918:data=8'h00;
14'h2919:data=8'h00;
14'h291a:data=8'h00;
14'h291b:data=8'h00;
14'h291c:data=8'h00;
14'h291d:data=8'h00;
14'h291e:data=8'h00;
14'h291f:data=8'h00;
14'h2920:data=8'h3E;
14'h2921:data=8'h00;
14'h2922:data=8'h00;
14'h2923:data=8'h00;
14'h2924:data=8'h00;
14'h2925:data=8'h00;
14'h2926:data=8'h78;
14'h2927:data=8'h00;
14'h2940:data=8'hFF;
14'h2941:data=8'hFF;
14'h2942:data=8'hFF;
14'h2943:data=8'hFF;
14'h2944:data=8'h80;
14'h2945:data=8'h00;
14'h2946:data=8'h00;
14'h2947:data=8'h00;
14'h2948:data=8'h00;
14'h2949:data=8'h00;
14'h294a:data=8'h03;
14'h294b:data=8'hFF;
14'h294c:data=8'hFF;
14'h294d:data=8'hFF;
14'h294e:data=8'hFF;
14'h294f:data=8'hFF;
14'h2950:data=8'hFF;
14'h2951:data=8'hFF;
14'h2952:data=8'hFF;
14'h2953:data=8'hFF;
14'h2954:data=8'h00;
14'h2955:data=8'h00;
14'h2956:data=8'h00;
14'h2957:data=8'h00;
14'h2958:data=8'h00;
14'h2959:data=8'h00;
14'h295a:data=8'h00;
14'h295b:data=8'h00;
14'h295c:data=8'h00;
14'h295d:data=8'h00;
14'h295e:data=8'h00;
14'h295f:data=8'h07;
14'h2960:data=8'hC0;
14'h2961:data=8'h00;
14'h2962:data=8'h00;
14'h2963:data=8'h00;
14'h2964:data=8'h00;
14'h2965:data=8'h03;
14'h2966:data=8'hC0;
14'h2967:data=8'h00;
14'h2980:data=8'hFF;
14'h2981:data=8'hFF;
14'h2982:data=8'hFF;
14'h2983:data=8'hFF;
14'h2984:data=8'h80;
14'h2985:data=8'h00;
14'h2986:data=8'h00;
14'h2987:data=8'h00;
14'h2988:data=8'h00;
14'h2989:data=8'h00;
14'h298a:data=8'h03;
14'h298b:data=8'hFF;
14'h298c:data=8'hFF;
14'h298d:data=8'hFF;
14'h298e:data=8'hFF;
14'h298f:data=8'hFF;
14'h2990:data=8'hFF;
14'h2991:data=8'hFF;
14'h2992:data=8'hFF;
14'h2993:data=8'hFF;
14'h2994:data=8'h00;
14'h2995:data=8'h00;
14'h2996:data=8'h00;
14'h2997:data=8'h00;
14'h2998:data=8'h00;
14'h2999:data=8'h00;
14'h299a:data=8'h00;
14'h299b:data=8'h00;
14'h299c:data=8'h00;
14'h299d:data=8'h00;
14'h299e:data=8'h01;
14'h299f:data=8'hF8;
14'h29a0:data=8'h00;
14'h29a1:data=8'h00;
14'h29a2:data=8'h00;
14'h29a3:data=8'h00;
14'h29a4:data=8'h00;
14'h29a5:data=8'h1C;
14'h29a6:data=8'h00;
14'h29a7:data=8'h00;
14'h29c0:data=8'hFF;
14'h29c1:data=8'hFF;
14'h29c2:data=8'hFF;
14'h29c3:data=8'hFF;
14'h29c4:data=8'h80;
14'h29c5:data=8'h00;
14'h29c6:data=8'h00;
14'h29c7:data=8'h00;
14'h29c8:data=8'h00;
14'h29c9:data=8'h00;
14'h29ca:data=8'h03;
14'h29cb:data=8'hFF;
14'h29cc:data=8'hFF;
14'h29cd:data=8'hFF;
14'h29ce:data=8'hFF;
14'h29cf:data=8'hFF;
14'h29d0:data=8'hFF;
14'h29d1:data=8'hFF;
14'h29d2:data=8'hFF;
14'h29d3:data=8'hFF;
14'h29d4:data=8'h00;
14'h29d5:data=8'h00;
14'h29d6:data=8'h00;
14'h29d7:data=8'h00;
14'h29d8:data=8'h00;
14'h29d9:data=8'h00;
14'h29da:data=8'h00;
14'h29db:data=8'h00;
14'h29dc:data=8'h00;
14'h29dd:data=8'h00;
14'h29de:data=8'h3F;
14'h29df:data=8'h00;
14'h29e0:data=8'h00;
14'h29e1:data=8'h00;
14'h29e2:data=8'h00;
14'h29e3:data=8'h00;
14'h29e4:data=8'h01;
14'h29e5:data=8'hE0;
14'h29e6:data=8'h00;
14'h29e7:data=8'h00;
14'h2a00:data=8'hFF;
14'h2a01:data=8'hFF;
14'h2a02:data=8'hFF;
14'h2a03:data=8'hFC;
14'h2a04:data=8'h00;
14'h2a05:data=8'h00;
14'h2a06:data=8'h00;
14'h2a07:data=8'h00;
14'h2a08:data=8'h00;
14'h2a09:data=8'h00;
14'h2a0a:data=8'h03;
14'h2a0b:data=8'hFF;
14'h2a0c:data=8'hFF;
14'h2a0d:data=8'hFF;
14'h2a0e:data=8'hFF;
14'h2a0f:data=8'hFF;
14'h2a10:data=8'hFF;
14'h2a11:data=8'hFF;
14'h2a12:data=8'hFF;
14'h2a13:data=8'hFF;
14'h2a14:data=8'h00;
14'h2a15:data=8'h00;
14'h2a16:data=8'h00;
14'h2a17:data=8'h00;
14'h2a18:data=8'h00;
14'h2a19:data=8'h00;
14'h2a1a:data=8'h00;
14'h2a1b:data=8'h00;
14'h2a1c:data=8'h00;
14'h2a1d:data=8'h07;
14'h2a1e:data=8'hE0;
14'h2a1f:data=8'h00;
14'h2a20:data=8'h00;
14'h2a21:data=8'h00;
14'h2a22:data=8'h00;
14'h2a23:data=8'h00;
14'h2a24:data=8'h0F;
14'h2a25:data=8'h00;
14'h2a26:data=8'h00;
14'h2a27:data=8'h00;
14'h2a40:data=8'hFF;
14'h2a41:data=8'hFF;
14'h2a42:data=8'hFF;
14'h2a43:data=8'hFC;
14'h2a44:data=8'h00;
14'h2a45:data=8'h00;
14'h2a46:data=8'h00;
14'h2a47:data=8'h00;
14'h2a48:data=8'h00;
14'h2a49:data=8'h00;
14'h2a4a:data=8'h03;
14'h2a4b:data=8'hFF;
14'h2a4c:data=8'hFF;
14'h2a4d:data=8'hFF;
14'h2a4e:data=8'hFF;
14'h2a4f:data=8'hFF;
14'h2a50:data=8'hFF;
14'h2a51:data=8'hFF;
14'h2a52:data=8'hFF;
14'h2a53:data=8'hFF;
14'h2a54:data=8'h00;
14'h2a55:data=8'h00;
14'h2a56:data=8'h00;
14'h2a57:data=8'h00;
14'h2a58:data=8'h00;
14'h2a59:data=8'h00;
14'h2a5a:data=8'h00;
14'h2a5b:data=8'h00;
14'h2a5c:data=8'h00;
14'h2a5d:data=8'hFC;
14'h2a5e:data=8'h00;
14'h2a5f:data=8'h00;
14'h2a60:data=8'h00;
14'h2a61:data=8'h00;
14'h2a62:data=8'h00;
14'h2a63:data=8'h00;
14'h2a64:data=8'h70;
14'h2a65:data=8'h00;
14'h2a66:data=8'h00;
14'h2a67:data=8'h00;
14'h2a80:data=8'hFF;
14'h2a81:data=8'hFF;
14'h2a82:data=8'hFF;
14'h2a83:data=8'hFC;
14'h2a84:data=8'h00;
14'h2a85:data=8'h00;
14'h2a86:data=8'h00;
14'h2a87:data=8'h00;
14'h2a88:data=8'h00;
14'h2a89:data=8'h00;
14'h2a8a:data=8'h03;
14'h2a8b:data=8'hFF;
14'h2a8c:data=8'hFF;
14'h2a8d:data=8'hFF;
14'h2a8e:data=8'hFF;
14'h2a8f:data=8'hFF;
14'h2a90:data=8'hFF;
14'h2a91:data=8'hFF;
14'h2a92:data=8'hFF;
14'h2a93:data=8'hFF;
14'h2a94:data=8'h00;
14'h2a95:data=8'h00;
14'h2a96:data=8'h00;
14'h2a97:data=8'h00;
14'h2a98:data=8'h00;
14'h2a99:data=8'h00;
14'h2a9a:data=8'h00;
14'h2a9b:data=8'h00;
14'h2a9c:data=8'h1F;
14'h2a9d:data=8'h00;
14'h2a9e:data=8'h00;
14'h2a9f:data=8'h00;
14'h2aa0:data=8'h00;
14'h2aa1:data=8'h00;
14'h2aa2:data=8'h00;
14'h2aa3:data=8'h03;
14'h2aa4:data=8'h80;
14'h2aa5:data=8'h00;
14'h2aa6:data=8'h00;
14'h2aa7:data=8'h00;
14'h2ac0:data=8'hFF;
14'h2ac1:data=8'hFF;
14'h2ac2:data=8'hFF;
14'h2ac3:data=8'hFC;
14'h2ac4:data=8'h00;
14'h2ac5:data=8'h00;
14'h2ac6:data=8'h00;
14'h2ac7:data=8'h00;
14'h2ac8:data=8'h00;
14'h2ac9:data=8'h00;
14'h2aca:data=8'h03;
14'h2acb:data=8'hFF;
14'h2acc:data=8'hFF;
14'h2acd:data=8'hFF;
14'h2ace:data=8'hFF;
14'h2acf:data=8'hFF;
14'h2ad0:data=8'hFF;
14'h2ad1:data=8'hFF;
14'h2ad2:data=8'hFF;
14'h2ad3:data=8'hFF;
14'h2ad4:data=8'h00;
14'h2ad5:data=8'h00;
14'h2ad6:data=8'h00;
14'h2ad7:data=8'h00;
14'h2ad8:data=8'h00;
14'h2ad9:data=8'h00;
14'h2ada:data=8'h00;
14'h2adb:data=8'h03;
14'h2adc:data=8'hE0;
14'h2add:data=8'h00;
14'h2ade:data=8'h00;
14'h2adf:data=8'h00;
14'h2ae0:data=8'h00;
14'h2ae1:data=8'h00;
14'h2ae2:data=8'h00;
14'h2ae3:data=8'h3C;
14'h2ae4:data=8'h00;
14'h2ae5:data=8'h00;
14'h2ae6:data=8'h00;
14'h2ae7:data=8'h00;
14'h2b00:data=8'hFF;
14'h2b01:data=8'hFF;
14'h2b02:data=8'hFF;
14'h2b03:data=8'hFC;
14'h2b04:data=8'h00;
14'h2b05:data=8'h00;
14'h2b06:data=8'h00;
14'h2b07:data=8'h00;
14'h2b08:data=8'h00;
14'h2b09:data=8'h00;
14'h2b0a:data=8'h03;
14'h2b0b:data=8'hFF;
14'h2b0c:data=8'hFF;
14'h2b0d:data=8'hFF;
14'h2b0e:data=8'hFF;
14'h2b0f:data=8'hFF;
14'h2b10:data=8'hFF;
14'h2b11:data=8'hFF;
14'h2b12:data=8'hFF;
14'h2b13:data=8'hF0;
14'h2b14:data=8'h00;
14'h2b15:data=8'h00;
14'h2b16:data=8'h00;
14'h2b17:data=8'h00;
14'h2b18:data=8'h00;
14'h2b19:data=8'h00;
14'h2b1a:data=8'h00;
14'h2b1b:data=8'hFC;
14'h2b1c:data=8'h00;
14'h2b1d:data=8'h00;
14'h2b1e:data=8'h00;
14'h2b1f:data=8'h00;
14'h2b20:data=8'h00;
14'h2b21:data=8'h00;
14'h2b22:data=8'h01;
14'h2b23:data=8'hE0;
14'h2b24:data=8'h00;
14'h2b25:data=8'h00;
14'h2b26:data=8'h00;
14'h2b27:data=8'h00;
14'h2b40:data=8'hFF;
14'h2b41:data=8'hFF;
14'h2b42:data=8'hFF;
14'h2b43:data=8'hFC;
14'h2b44:data=8'h00;
14'h2b45:data=8'h00;
14'h2b46:data=8'h00;
14'h2b47:data=8'h00;
14'h2b48:data=8'h00;
14'h2b49:data=8'h00;
14'h2b4a:data=8'h03;
14'h2b4b:data=8'hFF;
14'h2b4c:data=8'hFF;
14'h2b4d:data=8'hFF;
14'h2b4e:data=8'hFF;
14'h2b4f:data=8'hFF;
14'h2b50:data=8'hFF;
14'h2b51:data=8'hFF;
14'h2b52:data=8'hE0;
14'h2b53:data=8'h00;
14'h2b54:data=8'h00;
14'h2b55:data=8'h00;
14'h2b56:data=8'h00;
14'h2b57:data=8'h00;
14'h2b58:data=8'h00;
14'h2b59:data=8'h00;
14'h2b5a:data=8'h1F;
14'h2b5b:data=8'h80;
14'h2b5c:data=8'h00;
14'h2b5d:data=8'h00;
14'h2b5e:data=8'h00;
14'h2b5f:data=8'h00;
14'h2b60:data=8'h00;
14'h2b61:data=8'h00;
14'h2b62:data=8'h0E;
14'h2b63:data=8'h00;
14'h2b64:data=8'h00;
14'h2b65:data=8'h00;
14'h2b66:data=8'h00;
14'h2b67:data=8'h00;
14'h2b80:data=8'hFF;
14'h2b81:data=8'hFF;
14'h2b82:data=8'hFF;
14'h2b83:data=8'hC0;
14'h2b84:data=8'h00;
14'h2b85:data=8'h00;
14'h2b86:data=8'h00;
14'h2b87:data=8'h00;
14'h2b88:data=8'h00;
14'h2b89:data=8'h00;
14'h2b8a:data=8'h03;
14'h2b8b:data=8'hFF;
14'h2b8c:data=8'hFF;
14'h2b8d:data=8'hFF;
14'h2b8e:data=8'hFF;
14'h2b8f:data=8'hFF;
14'h2b90:data=8'hFF;
14'h2b91:data=8'hC0;
14'h2b92:data=8'h00;
14'h2b93:data=8'h00;
14'h2b94:data=8'h00;
14'h2b95:data=8'h00;
14'h2b96:data=8'h00;
14'h2b97:data=8'h00;
14'h2b98:data=8'h00;
14'h2b99:data=8'h03;
14'h2b9a:data=8'hF0;
14'h2b9b:data=8'h00;
14'h2b9c:data=8'h00;
14'h2b9d:data=8'h00;
14'h2b9e:data=8'h00;
14'h2b9f:data=8'h00;
14'h2ba0:data=8'h00;
14'h2ba1:data=8'h00;
14'h2ba2:data=8'hF0;
14'h2ba3:data=8'h00;
14'h2ba4:data=8'h00;
14'h2ba5:data=8'h00;
14'h2ba6:data=8'h00;
14'h2ba7:data=8'h00;
14'h2bc0:data=8'hFF;
14'h2bc1:data=8'hFF;
14'h2bc2:data=8'hFF;
14'h2bc3:data=8'h80;
14'h2bc4:data=8'h00;
14'h2bc5:data=8'h00;
14'h2bc6:data=8'h00;
14'h2bc7:data=8'h00;
14'h2bc8:data=8'h00;
14'h2bc9:data=8'h00;
14'h2bca:data=8'h03;
14'h2bcb:data=8'hFF;
14'h2bcc:data=8'hFF;
14'h2bcd:data=8'hFF;
14'h2bce:data=8'hFF;
14'h2bcf:data=8'hFF;
14'h2bd0:data=8'h80;
14'h2bd1:data=8'h00;
14'h2bd2:data=8'h00;
14'h2bd3:data=8'h00;
14'h2bd4:data=8'h00;
14'h2bd5:data=8'h00;
14'h2bd6:data=8'h00;
14'h2bd7:data=8'h00;
14'h2bd8:data=8'h00;
14'h2bd9:data=8'h7C;
14'h2bda:data=8'h00;
14'h2bdb:data=8'h00;
14'h2bdc:data=8'h00;
14'h2bdd:data=8'h00;
14'h2bde:data=8'h00;
14'h2bdf:data=8'h00;
14'h2be0:data=8'h00;
14'h2be1:data=8'h07;
14'h2be2:data=8'h80;
14'h2be3:data=8'h00;
14'h2be4:data=8'h00;
14'h2be5:data=8'h00;
14'h2be6:data=8'h00;
14'h2be7:data=8'h00;
14'h2c00:data=8'hFF;
14'h2c01:data=8'hFF;
14'h2c02:data=8'hFF;
14'h2c03:data=8'h80;
14'h2c04:data=8'h00;
14'h2c05:data=8'h00;
14'h2c06:data=8'h00;
14'h2c07:data=8'h00;
14'h2c08:data=8'h00;
14'h2c09:data=8'h00;
14'h2c0a:data=8'h03;
14'h2c0b:data=8'hFF;
14'h2c0c:data=8'hFF;
14'h2c0d:data=8'hFF;
14'h2c0e:data=8'hFF;
14'h2c0f:data=8'h00;
14'h2c10:data=8'h00;
14'h2c11:data=8'h00;
14'h2c12:data=8'h00;
14'h2c13:data=8'h00;
14'h2c14:data=8'h00;
14'h2c15:data=8'h00;
14'h2c16:data=8'h00;
14'h2c17:data=8'h00;
14'h2c18:data=8'h0F;
14'h2c19:data=8'h80;
14'h2c1a:data=8'h00;
14'h2c1b:data=8'h00;
14'h2c1c:data=8'h00;
14'h2c1d:data=8'h00;
14'h2c1e:data=8'h00;
14'h2c1f:data=8'h00;
14'h2c20:data=8'h00;
14'h2c21:data=8'h38;
14'h2c22:data=8'h00;
14'h2c23:data=8'h00;
14'h2c24:data=8'h00;
14'h2c25:data=8'h00;
14'h2c26:data=8'h00;
14'h2c27:data=8'h00;
14'h2c40:data=8'hFF;
14'h2c41:data=8'hFF;
14'h2c42:data=8'hFF;
14'h2c43:data=8'h80;
14'h2c44:data=8'h00;
14'h2c45:data=8'h00;
14'h2c46:data=8'h00;
14'h2c47:data=8'h00;
14'h2c48:data=8'h00;
14'h2c49:data=8'h00;
14'h2c4a:data=8'h00;
14'h2c4b:data=8'h1F;
14'h2c4c:data=8'hFF;
14'h2c4d:data=8'hFE;
14'h2c4e:data=8'h00;
14'h2c4f:data=8'h00;
14'h2c50:data=8'h00;
14'h2c51:data=8'h00;
14'h2c52:data=8'h00;
14'h2c53:data=8'h00;
14'h2c54:data=8'h00;
14'h2c55:data=8'h00;
14'h2c56:data=8'h00;
14'h2c57:data=8'h03;
14'h2c58:data=8'hF0;
14'h2c59:data=8'h00;
14'h2c5a:data=8'h00;
14'h2c5b:data=8'h00;
14'h2c5c:data=8'h00;
14'h2c5d:data=8'h00;
14'h2c5e:data=8'h00;
14'h2c5f:data=8'h00;
14'h2c60:data=8'h03;
14'h2c61:data=8'hC0;
14'h2c62:data=8'h00;
14'h2c63:data=8'h00;
14'h2c64:data=8'h00;
14'h2c65:data=8'h00;
14'h2c66:data=8'h00;
14'h2c67:data=8'h00;
14'h2c80:data=8'hFF;
14'h2c81:data=8'hFF;
14'h2c82:data=8'hFF;
14'h2c83:data=8'h80;
14'h2c84:data=8'h00;
14'h2c85:data=8'h00;
14'h2c86:data=8'h00;
14'h2c87:data=8'h00;
14'h2c88:data=8'h00;
14'h2c89:data=8'h00;
14'h2c8a:data=8'h00;
14'h2c8b:data=8'h1F;
14'h2c8c:data=8'hFC;
14'h2c8d:data=8'h00;
14'h2c8e:data=8'h00;
14'h2c8f:data=8'h00;
14'h2c90:data=8'h00;
14'h2c91:data=8'h00;
14'h2c92:data=8'h00;
14'h2c93:data=8'h00;
14'h2c94:data=8'h00;
14'h2c95:data=8'h00;
14'h2c96:data=8'h00;
14'h2c97:data=8'h7E;
14'h2c98:data=8'h00;
14'h2c99:data=8'h00;
14'h2c9a:data=8'h00;
14'h2c9b:data=8'h00;
14'h2c9c:data=8'h00;
14'h2c9d:data=8'h00;
14'h2c9e:data=8'h00;
14'h2c9f:data=8'h00;
14'h2ca0:data=8'h7E;
14'h2ca1:data=8'h00;
14'h2ca2:data=8'h00;
14'h2ca3:data=8'h00;
14'h2ca4:data=8'h00;
14'h2ca5:data=8'h00;
14'h2ca6:data=8'h00;
14'h2ca7:data=8'h00;
14'h2cc0:data=8'h00;
14'h2cc1:data=8'h00;
14'h2cc2:data=8'h00;
14'h2cc3:data=8'h00;
14'h2cc4:data=8'h00;
14'h2cc5:data=8'h00;
14'h2cc6:data=8'h00;
14'h2cc7:data=8'h00;
14'h2cc8:data=8'h00;
14'h2cc9:data=8'h00;
14'h2cca:data=8'h00;
14'h2ccb:data=8'h08;
14'h2ccc:data=8'h00;
14'h2ccd:data=8'h00;
14'h2cce:data=8'h00;
14'h2ccf:data=8'h00;
14'h2cd0:data=8'h00;
14'h2cd1:data=8'h00;
14'h2cd2:data=8'h00;
14'h2cd3:data=8'h00;
14'h2cd4:data=8'h00;
14'h2cd5:data=8'h00;
14'h2cd6:data=8'h0F;
14'h2cd7:data=8'hC0;
14'h2cd8:data=8'h00;
14'h2cd9:data=8'h00;
14'h2cda:data=8'h00;
14'h2cdb:data=8'h00;
14'h2cdc:data=8'h00;
14'h2cdd:data=8'h00;
14'h2cde:data=8'h00;
14'h2cdf:data=8'h0F;
14'h2ce0:data=8'hC0;
14'h2ce1:data=8'h00;
14'h2ce2:data=8'h00;
14'h2ce3:data=8'h00;
14'h2ce4:data=8'h00;
14'h2ce5:data=8'h00;
14'h2ce6:data=8'h00;
14'h2ce7:data=8'h00;
14'h2d00:data=8'h00;
14'h2d01:data=8'h00;
14'h2d02:data=8'h00;
14'h2d03:data=8'h00;
14'h2d04:data=8'h00;
14'h2d05:data=8'h00;
14'h2d06:data=8'h00;
14'h2d07:data=8'h00;
14'h2d08:data=8'h00;
14'h2d09:data=8'h00;
14'h2d0a:data=8'h00;
14'h2d0b:data=8'h00;
14'h2d0c:data=8'h00;
14'h2d0d:data=8'h00;
14'h2d0e:data=8'h00;
14'h2d0f:data=8'h00;
14'h2d10:data=8'h00;
14'h2d11:data=8'h00;
14'h2d12:data=8'h00;
14'h2d13:data=8'h00;
14'h2d14:data=8'h00;
14'h2d15:data=8'h01;
14'h2d16:data=8'hF8;
14'h2d17:data=8'h00;
14'h2d18:data=8'h00;
14'h2d19:data=8'h00;
14'h2d1a:data=8'h00;
14'h2d1b:data=8'h00;
14'h2d1c:data=8'h00;
14'h2d1d:data=8'h00;
14'h2d1e:data=8'h01;
14'h2d1f:data=8'hF8;
14'h2d20:data=8'h00;
14'h2d21:data=8'h00;
14'h2d22:data=8'h00;
14'h2d23:data=8'h00;
14'h2d24:data=8'h00;
14'h2d25:data=8'h00;
14'h2d26:data=8'h00;
14'h2d27:data=8'h00;
14'h2d40:data=8'h00;
14'h2d41:data=8'h00;
14'h2d42:data=8'h00;
14'h2d43:data=8'h00;
14'h2d44:data=8'h00;
14'h2d45:data=8'h00;
14'h2d46:data=8'h00;
14'h2d47:data=8'h00;
14'h2d48:data=8'h00;
14'h2d49:data=8'h00;
14'h2d4a:data=8'h00;
14'h2d4b:data=8'h00;
14'h2d4c:data=8'h00;
14'h2d4d:data=8'h00;
14'h2d4e:data=8'h00;
14'h2d4f:data=8'h00;
14'h2d50:data=8'h00;
14'h2d51:data=8'h00;
14'h2d52:data=8'h00;
14'h2d53:data=8'h00;
14'h2d54:data=8'h00;
14'h2d55:data=8'h3C;
14'h2d56:data=8'h00;
14'h2d57:data=8'h00;
14'h2d58:data=8'h00;
14'h2d59:data=8'h00;
14'h2d5a:data=8'h00;
14'h2d5b:data=8'h00;
14'h2d5c:data=8'h00;
14'h2d5d:data=8'h00;
14'h2d5e:data=8'h3C;
14'h2d5f:data=8'h00;
14'h2d60:data=8'h00;
14'h2d61:data=8'h00;
14'h2d62:data=8'h00;
14'h2d63:data=8'h00;
14'h2d64:data=8'h00;
14'h2d65:data=8'h00;
14'h2d66:data=8'h00;
14'h2d67:data=8'h00;
14'h2d80:data=8'h00;
14'h2d81:data=8'h00;
14'h2d82:data=8'h00;
14'h2d83:data=8'h00;
14'h2d84:data=8'h00;
14'h2d85:data=8'h00;
14'h2d86:data=8'h00;
14'h2d87:data=8'h00;
14'h2d88:data=8'h00;
14'h2d89:data=8'h00;
14'h2d8a:data=8'h00;
14'h2d8b:data=8'h00;
14'h2d8c:data=8'h00;
14'h2d8d:data=8'h00;
14'h2d8e:data=8'h00;
14'h2d8f:data=8'h00;
14'h2d90:data=8'h00;
14'h2d91:data=8'h00;
14'h2d92:data=8'h00;
14'h2d93:data=8'h00;
14'h2d94:data=8'h07;
14'h2d95:data=8'h80;
14'h2d96:data=8'h00;
14'h2d97:data=8'h00;
14'h2d98:data=8'h00;
14'h2d99:data=8'h00;
14'h2d9a:data=8'h00;
14'h2d9b:data=8'h00;
14'h2d9c:data=8'h00;
14'h2d9d:data=8'h07;
14'h2d9e:data=8'h80;
14'h2d9f:data=8'h00;
14'h2da0:data=8'h00;
14'h2da1:data=8'h00;
14'h2da2:data=8'h00;
14'h2da3:data=8'h00;
14'h2da4:data=8'h00;
14'h2da5:data=8'h00;
14'h2da6:data=8'h00;
14'h2da7:data=8'h00;
14'h2dc0:data=8'h00;
14'h2dc1:data=8'h00;
14'h2dc2:data=8'h00;
14'h2dc3:data=8'h00;
14'h2dc4:data=8'h00;
14'h2dc5:data=8'h00;
14'h2dc6:data=8'h00;
14'h2dc7:data=8'h00;
14'h2dc8:data=8'h00;
14'h2dc9:data=8'h00;
14'h2dca:data=8'h00;
14'h2dcb:data=8'h00;
14'h2dcc:data=8'h00;
14'h2dcd:data=8'h00;
14'h2dce:data=8'h00;
14'h2dcf:data=8'h00;
14'h2dd0:data=8'h00;
14'h2dd1:data=8'h00;
14'h2dd2:data=8'h00;
14'h2dd3:data=8'h01;
14'h2dd4:data=8'hF0;
14'h2dd5:data=8'h00;
14'h2dd6:data=8'h00;
14'h2dd7:data=8'h00;
14'h2dd8:data=8'h00;
14'h2dd9:data=8'h00;
14'h2dda:data=8'h00;
14'h2ddb:data=8'h00;
14'h2ddc:data=8'h00;
14'h2ddd:data=8'hF0;
14'h2dde:data=8'h00;
14'h2ddf:data=8'h00;
14'h2de0:data=8'h00;
14'h2de1:data=8'h00;
14'h2de2:data=8'h00;
14'h2de3:data=8'h00;
14'h2de4:data=8'h00;
14'h2de5:data=8'h00;
14'h2de6:data=8'h00;
14'h2de7:data=8'h00;
14'h2e00:data=8'h00;
14'h2e01:data=8'h00;
14'h2e02:data=8'h00;
14'h2e03:data=8'h00;
14'h2e04:data=8'h00;
14'h2e05:data=8'h00;
14'h2e06:data=8'h00;
14'h2e07:data=8'h00;
14'h2e08:data=8'h00;
14'h2e09:data=8'h00;
14'h2e0a:data=8'h00;
14'h2e0b:data=8'h00;
14'h2e0c:data=8'h00;
14'h2e0d:data=8'h00;
14'h2e0e:data=8'h00;
14'h2e0f:data=8'h00;
14'h2e10:data=8'h00;
14'h2e11:data=8'h00;
14'h2e12:data=8'h00;
14'h2e13:data=8'h3C;
14'h2e14:data=8'h00;
14'h2e15:data=8'h00;
14'h2e16:data=8'h00;
14'h2e17:data=8'h00;
14'h2e18:data=8'h00;
14'h2e19:data=8'h00;
14'h2e1a:data=8'h00;
14'h2e1b:data=8'h00;
14'h2e1c:data=8'h1E;
14'h2e1d:data=8'h00;
14'h2e1e:data=8'h00;
14'h2e1f:data=8'h00;
14'h2e20:data=8'h00;
14'h2e21:data=8'h00;
14'h2e22:data=8'h00;
14'h2e23:data=8'h00;
14'h2e24:data=8'h00;
14'h2e25:data=8'h00;
14'h2e26:data=8'h00;
14'h2e27:data=8'h00;
14'h2e40:data=8'h00;
14'h2e41:data=8'h00;
14'h2e42:data=8'h00;
14'h2e43:data=8'h00;
14'h2e44:data=8'h00;
14'h2e45:data=8'h00;
14'h2e46:data=8'h00;
14'h2e47:data=8'h00;
14'h2e48:data=8'h00;
14'h2e49:data=8'h00;
14'h2e4a:data=8'h00;
14'h2e4b:data=8'h00;
14'h2e4c:data=8'h00;
14'h2e4d:data=8'h00;
14'h2e4e:data=8'h00;
14'h2e4f:data=8'h00;
14'h2e50:data=8'h00;
14'h2e51:data=8'h00;
14'h2e52:data=8'h07;
14'h2e53:data=8'h80;
14'h2e54:data=8'h00;
14'h2e55:data=8'h00;
14'h2e56:data=8'h00;
14'h2e57:data=8'h00;
14'h2e58:data=8'h00;
14'h2e59:data=8'h00;
14'h2e5a:data=8'h00;
14'h2e5b:data=8'h03;
14'h2e5c:data=8'hC0;
14'h2e5d:data=8'h00;
14'h2e5e:data=8'h00;
14'h2e5f:data=8'h00;
14'h2e60:data=8'h00;
14'h2e61:data=8'h00;
14'h2e62:data=8'h00;
14'h2e63:data=8'h00;
14'h2e64:data=8'h00;
14'h2e65:data=8'h00;
14'h2e66:data=8'h00;
14'h2e67:data=8'h00;
14'h2e80:data=8'h00;
14'h2e81:data=8'h00;
14'h2e82:data=8'h00;
14'h2e83:data=8'h00;
14'h2e84:data=8'h00;
14'h2e85:data=8'h00;
14'h2e86:data=8'h00;
14'h2e87:data=8'h00;
14'h2e88:data=8'h00;
14'h2e89:data=8'h00;
14'h2e8a:data=8'h00;
14'h2e8b:data=8'h00;
14'h2e8c:data=8'h00;
14'h2e8d:data=8'h00;
14'h2e8e:data=8'h00;
14'h2e8f:data=8'h00;
14'h2e90:data=8'h00;
14'h2e91:data=8'h00;
14'h2e92:data=8'hF0;
14'h2e93:data=8'h00;
14'h2e94:data=8'h00;
14'h2e95:data=8'h00;
14'h2e96:data=8'h00;
14'h2e97:data=8'h00;
14'h2e98:data=8'h00;
14'h2e99:data=8'h00;
14'h2e9a:data=8'h00;
14'h2e9b:data=8'h78;
14'h2e9c:data=8'h00;
14'h2e9d:data=8'h00;
14'h2e9e:data=8'h00;
14'h2e9f:data=8'h00;
14'h2ea0:data=8'h00;
14'h2ea1:data=8'h00;
14'h2ea2:data=8'h00;
14'h2ea3:data=8'h00;
14'h2ea4:data=8'h00;
14'h2ea5:data=8'h00;
14'h2ea6:data=8'h00;
14'h2ea7:data=8'h00;
14'h2ec0:data=8'h00;
14'h2ec1:data=8'h00;
14'h2ec2:data=8'h00;
14'h2ec3:data=8'h00;
14'h2ec4:data=8'h00;
14'h2ec5:data=8'h00;
14'h2ec6:data=8'h00;
14'h2ec7:data=8'h00;
14'h2ec8:data=8'h00;
14'h2ec9:data=8'h00;
14'h2eca:data=8'h00;
14'h2ecb:data=8'h00;
14'h2ecc:data=8'h00;
14'h2ecd:data=8'h00;
14'h2ece:data=8'h00;
14'h2ecf:data=8'h00;
14'h2ed0:data=8'h00;
14'h2ed1:data=8'h1E;
14'h2ed2:data=8'h00;
14'h2ed3:data=8'h00;
14'h2ed4:data=8'h00;
14'h2ed5:data=8'h00;
14'h2ed6:data=8'h00;
14'h2ed7:data=8'h00;
14'h2ed8:data=8'h00;
14'h2ed9:data=8'h00;
14'h2eda:data=8'h0F;
14'h2edb:data=8'h00;
14'h2edc:data=8'h00;
14'h2edd:data=8'h00;
14'h2ede:data=8'h00;
14'h2edf:data=8'h00;
14'h2ee0:data=8'h00;
14'h2ee1:data=8'h00;
14'h2ee2:data=8'h00;
14'h2ee3:data=8'h00;
14'h2ee4:data=8'h00;
14'h2ee5:data=8'h00;
14'h2ee6:data=8'h00;
14'h2ee7:data=8'h00;
14'h2f00:data=8'h00;
14'h2f01:data=8'h00;
14'h2f02:data=8'h00;
14'h2f03:data=8'h00;
14'h2f04:data=8'h00;
14'h2f05:data=8'h00;
14'h2f06:data=8'h00;
14'h2f07:data=8'h00;
14'h2f08:data=8'h00;
14'h2f09:data=8'h00;
14'h2f0a:data=8'h00;
14'h2f0b:data=8'h00;
14'h2f0c:data=8'h00;
14'h2f0d:data=8'h00;
14'h2f0e:data=8'h00;
14'h2f0f:data=8'h00;
14'h2f10:data=8'h03;
14'h2f11:data=8'h80;
14'h2f12:data=8'h00;
14'h2f13:data=8'h00;
14'h2f14:data=8'h00;
14'h2f15:data=8'h00;
14'h2f16:data=8'h00;
14'h2f17:data=8'h00;
14'h2f18:data=8'h00;
14'h2f19:data=8'h01;
14'h2f1a:data=8'hE0;
14'h2f1b:data=8'h00;
14'h2f1c:data=8'h00;
14'h2f1d:data=8'h00;
14'h2f1e:data=8'h00;
14'h2f1f:data=8'h00;
14'h2f20:data=8'h00;
14'h2f21:data=8'h00;
14'h2f22:data=8'h00;
14'h2f23:data=8'h00;
14'h2f24:data=8'h00;
14'h2f25:data=8'h00;
14'h2f26:data=8'h00;
14'h2f27:data=8'h00;
14'h2f40:data=8'h00;
14'h2f41:data=8'h00;
14'h2f42:data=8'h00;
14'h2f43:data=8'h00;
14'h2f44:data=8'h00;
14'h2f45:data=8'h00;
14'h2f46:data=8'h00;
14'h2f47:data=8'h00;
14'h2f48:data=8'h00;
14'h2f49:data=8'h00;
14'h2f4a:data=8'h00;
14'h2f4b:data=8'h00;
14'h2f4c:data=8'h00;
14'h2f4d:data=8'h00;
14'h2f4e:data=8'h00;
14'h2f4f:data=8'h00;
14'h2f50:data=8'hF8;
14'h2f51:data=8'h00;
14'h2f52:data=8'h00;
14'h2f53:data=8'h00;
14'h2f54:data=8'h00;
14'h2f55:data=8'h00;
14'h2f56:data=8'h00;
14'h2f57:data=8'h00;
14'h2f58:data=8'h00;
14'h2f59:data=8'h3C;
14'h2f5a:data=8'h00;
14'h2f5b:data=8'h00;
14'h2f5c:data=8'h00;
14'h2f5d:data=8'h00;
14'h2f5e:data=8'h00;
14'h2f5f:data=8'h00;
14'h2f60:data=8'h00;
14'h2f61:data=8'h00;
14'h2f62:data=8'h00;
14'h2f63:data=8'h00;
14'h2f64:data=8'h00;
14'h2f65:data=8'h00;
14'h2f66:data=8'h00;
14'h2f67:data=8'h00;
14'h2f80:data=8'h00;
14'h2f81:data=8'h00;
14'h2f82:data=8'h00;
14'h2f83:data=8'h00;
14'h2f84:data=8'h00;
14'h2f85:data=8'h00;
14'h2f86:data=8'h00;
14'h2f87:data=8'h00;
14'h2f88:data=8'h00;
14'h2f89:data=8'h00;
14'h2f8a:data=8'h00;
14'h2f8b:data=8'h00;
14'h2f8c:data=8'h00;
14'h2f8d:data=8'h00;
14'h2f8e:data=8'h00;
14'h2f8f:data=8'h3E;
14'h2f90:data=8'h00;
14'h2f91:data=8'h00;
14'h2f92:data=8'h00;
14'h2f93:data=8'h00;
14'h2f94:data=8'h00;
14'h2f95:data=8'h00;
14'h2f96:data=8'h00;
14'h2f97:data=8'h00;
14'h2f98:data=8'h1F;
14'h2f99:data=8'h80;
14'h2f9a:data=8'h00;
14'h2f9b:data=8'h00;
14'h2f9c:data=8'h00;
14'h2f9d:data=8'h00;
14'h2f9e:data=8'h00;
14'h2f9f:data=8'h00;
14'h2fa0:data=8'h00;
14'h2fa1:data=8'h00;
14'h2fa2:data=8'h00;
14'h2fa3:data=8'h00;
14'h2fa4:data=8'h00;
14'h2fa5:data=8'h00;
14'h2fa6:data=8'h00;
14'h2fa7:data=8'h00;
14'h2fc0:data=8'h00;
14'h2fc1:data=8'h00;
14'h2fc2:data=8'h00;
14'h2fc3:data=8'h00;
14'h2fc4:data=8'h00;
14'h2fc5:data=8'h00;
14'h2fc6:data=8'h00;
14'h2fc7:data=8'h00;
14'h2fc8:data=8'h00;
14'h2fc9:data=8'h00;
14'h2fca:data=8'h00;
14'h2fcb:data=8'h00;
14'h2fcc:data=8'h00;
14'h2fcd:data=8'h00;
14'h2fce:data=8'h07;
14'h2fcf:data=8'hC0;
14'h2fd0:data=8'h00;
14'h2fd1:data=8'h00;
14'h2fd2:data=8'h00;
14'h2fd3:data=8'h00;
14'h2fd4:data=8'h00;
14'h2fd5:data=8'h00;
14'h2fd6:data=8'h00;
14'h2fd7:data=8'h03;
14'h2fd8:data=8'hF0;
14'h2fd9:data=8'h00;
14'h2fda:data=8'h00;
14'h2fdb:data=8'h00;
14'h2fdc:data=8'h00;
14'h2fdd:data=8'h00;
14'h2fde:data=8'h00;
14'h2fdf:data=8'h00;
14'h2fe0:data=8'h00;
14'h2fe1:data=8'h00;
14'h2fe2:data=8'h00;
14'h2fe3:data=8'h00;
14'h2fe4:data=8'h00;
14'h2fe5:data=8'h00;
14'h2fe6:data=8'h00;
14'h2fe7:data=8'h00;
14'h3000:data=8'h00;
14'h3001:data=8'h00;
14'h3002:data=8'h00;
14'h3003:data=8'h00;
14'h3004:data=8'h00;
14'h3005:data=8'h00;
14'h3006:data=8'h00;
14'h3007:data=8'h00;
14'h3008:data=8'h00;
14'h3009:data=8'h00;
14'h300a:data=8'h00;
14'h300b:data=8'h00;
14'h300c:data=8'h00;
14'h300d:data=8'h00;
14'h300e:data=8'hF8;
14'h300f:data=8'h00;
14'h3010:data=8'h00;
14'h3011:data=8'h00;
14'h3012:data=8'h00;
14'h3013:data=8'h00;
14'h3014:data=8'h00;
14'h3015:data=8'h00;
14'h3016:data=8'h00;
14'h3017:data=8'h7E;
14'h3018:data=8'h00;
14'h3019:data=8'h00;
14'h301a:data=8'h00;
14'h301b:data=8'h00;
14'h301c:data=8'h00;
14'h301d:data=8'h00;
14'h301e:data=8'h00;
14'h301f:data=8'h00;
14'h3020:data=8'h00;
14'h3021:data=8'h00;
14'h3022:data=8'h00;
14'h3023:data=8'h00;
14'h3024:data=8'h00;
14'h3025:data=8'h00;
14'h3026:data=8'h00;
14'h3027:data=8'h00;
14'h3040:data=8'h00;
14'h3041:data=8'h00;
14'h3042:data=8'h00;
14'h3043:data=8'h00;
14'h3044:data=8'h00;
14'h3045:data=8'h00;
14'h3046:data=8'h00;
14'h3047:data=8'h00;
14'h3048:data=8'h00;
14'h3049:data=8'h00;
14'h304a:data=8'h00;
14'h304b:data=8'h00;
14'h304c:data=8'h00;
14'h304d:data=8'h1F;
14'h304e:data=8'h80;
14'h304f:data=8'h00;
14'h3050:data=8'h00;
14'h3051:data=8'h00;
14'h3052:data=8'h00;
14'h3053:data=8'h00;
14'h3054:data=8'h00;
14'h3055:data=8'h00;
14'h3056:data=8'h0F;
14'h3057:data=8'hC0;
14'h3058:data=8'h00;
14'h3059:data=8'h00;
14'h305a:data=8'h00;
14'h305b:data=8'h00;
14'h305c:data=8'h00;
14'h305d:data=8'h00;
14'h305e:data=8'h00;
14'h305f:data=8'h00;
14'h3060:data=8'h00;
14'h3061:data=8'h00;
14'h3062:data=8'h00;
14'h3063:data=8'h00;
14'h3064:data=8'h00;
14'h3065:data=8'h00;
14'h3066:data=8'h00;
14'h3067:data=8'h00;
14'h3080:data=8'h00;
14'h3081:data=8'h00;
14'h3082:data=8'h00;
14'h3083:data=8'h00;
14'h3084:data=8'h00;
14'h3085:data=8'h00;
14'h3086:data=8'h00;
14'h3087:data=8'h00;
14'h3088:data=8'h00;
14'h3089:data=8'h00;
14'h308a:data=8'h00;
14'h308b:data=8'h00;
14'h308c:data=8'h03;
14'h308d:data=8'hE0;
14'h308e:data=8'h00;
14'h308f:data=8'h00;
14'h3090:data=8'h00;
14'h3091:data=8'h00;
14'h3092:data=8'h00;
14'h3093:data=8'h00;
14'h3094:data=8'h00;
14'h3095:data=8'h01;
14'h3096:data=8'hF8;
14'h3097:data=8'h00;
14'h3098:data=8'h00;
14'h3099:data=8'h00;
14'h309a:data=8'h00;
14'h309b:data=8'h00;
14'h309c:data=8'h00;
14'h309d:data=8'h00;
14'h309e:data=8'h00;
14'h309f:data=8'h00;
14'h30a0:data=8'h00;
14'h30a1:data=8'h00;
14'h30a2:data=8'h00;
14'h30a3:data=8'h00;
14'h30a4:data=8'h00;
14'h30a5:data=8'h00;
14'h30a6:data=8'h00;
14'h30a7:data=8'h00;
14'h30c0:data=8'h00;
14'h30c1:data=8'h00;
14'h30c2:data=8'h00;
14'h30c3:data=8'h00;
14'h30c4:data=8'h00;
14'h30c5:data=8'h00;
14'h30c6:data=8'h00;
14'h30c7:data=8'h00;
14'h30c8:data=8'h00;
14'h30c9:data=8'h00;
14'h30ca:data=8'h00;
14'h30cb:data=8'h00;
14'h30cc:data=8'h7C;
14'h30cd:data=8'h00;
14'h30ce:data=8'h00;
14'h30cf:data=8'h00;
14'h30d0:data=8'h00;
14'h30d1:data=8'h00;
14'h30d2:data=8'h00;
14'h30d3:data=8'h00;
14'h30d4:data=8'h00;
14'h30d5:data=8'h3E;
14'h30d6:data=8'h00;
14'h30d7:data=8'h00;
14'h30d8:data=8'h00;
14'h30d9:data=8'h00;
14'h30da:data=8'h00;
14'h30db:data=8'h00;
14'h30dc:data=8'h00;
14'h30dd:data=8'h00;
14'h30de:data=8'h00;
14'h30df:data=8'h00;
14'h30e0:data=8'h00;
14'h30e1:data=8'h00;
14'h30e2:data=8'h00;
14'h30e3:data=8'h00;
14'h30e4:data=8'h00;
14'h30e5:data=8'h00;
14'h30e6:data=8'h00;
14'h30e7:data=8'h00;
14'h3100:data=8'h00;
14'h3101:data=8'h00;
14'h3102:data=8'h00;
14'h3103:data=8'h00;
14'h3104:data=8'h00;
14'h3105:data=8'h00;
14'h3106:data=8'h00;
14'h3107:data=8'h00;
14'h3108:data=8'h00;
14'h3109:data=8'h00;
14'h310a:data=8'h00;
14'h310b:data=8'h0F;
14'h310c:data=8'h80;
14'h310d:data=8'h00;
14'h310e:data=8'h00;
14'h310f:data=8'h00;
14'h3110:data=8'h00;
14'h3111:data=8'h00;
14'h3112:data=8'h00;
14'h3113:data=8'h00;
14'h3114:data=8'h07;
14'h3115:data=8'hC0;
14'h3116:data=8'h00;
14'h3117:data=8'h00;
14'h3118:data=8'h00;
14'h3119:data=8'h00;
14'h311a:data=8'h00;
14'h311b:data=8'h00;
14'h311c:data=8'h00;
14'h311d:data=8'h00;
14'h311e:data=8'h00;
14'h311f:data=8'h00;
14'h3120:data=8'h00;
14'h3121:data=8'h00;
14'h3122:data=8'h00;
14'h3123:data=8'h00;
14'h3124:data=8'h00;
14'h3125:data=8'h00;
14'h3126:data=8'h00;
14'h3127:data=8'h00;
14'h3140:data=8'h00;
14'h3141:data=8'h00;
14'h3142:data=8'h00;
14'h3143:data=8'h00;
14'h3144:data=8'h00;
14'h3145:data=8'h00;
14'h3146:data=8'h00;
14'h3147:data=8'h00;
14'h3148:data=8'h00;
14'h3149:data=8'h00;
14'h314a:data=8'h01;
14'h314b:data=8'hF8;
14'h314c:data=8'h00;
14'h314d:data=8'h00;
14'h314e:data=8'h00;
14'h314f:data=8'h00;
14'h3150:data=8'h00;
14'h3151:data=8'h00;
14'h3152:data=8'h00;
14'h3153:data=8'h00;
14'h3154:data=8'hFC;
14'h3155:data=8'h00;
14'h3156:data=8'h00;
14'h3157:data=8'h00;
14'h3158:data=8'h00;
14'h3159:data=8'h00;
14'h315a:data=8'h00;
14'h315b:data=8'h00;
14'h315c:data=8'h00;
14'h315d:data=8'h00;
14'h315e:data=8'h00;
14'h315f:data=8'h00;
14'h3160:data=8'h00;
14'h3161:data=8'h00;
14'h3162:data=8'h00;
14'h3163:data=8'h00;
14'h3164:data=8'h00;
14'h3165:data=8'h00;
14'h3166:data=8'h00;
14'h3167:data=8'h00;
14'h3180:data=8'h00;
14'h3181:data=8'h00;
14'h3182:data=8'h00;
14'h3183:data=8'h00;
14'h3184:data=8'h00;
14'h3185:data=8'h00;
14'h3186:data=8'h00;
14'h3187:data=8'h00;
14'h3188:data=8'h00;
14'h3189:data=8'h00;
14'h318a:data=8'h3E;
14'h318b:data=8'h00;
14'h318c:data=8'h00;
14'h318d:data=8'h00;
14'h318e:data=8'h00;
14'h318f:data=8'h00;
14'h3190:data=8'h00;
14'h3191:data=8'h00;
14'h3192:data=8'h00;
14'h3193:data=8'h1F;
14'h3194:data=8'h00;
14'h3195:data=8'h00;
14'h3196:data=8'h00;
14'h3197:data=8'h00;
14'h3198:data=8'h00;
14'h3199:data=8'h00;
14'h319a:data=8'h00;
14'h319b:data=8'h00;
14'h319c:data=8'h00;
14'h319d:data=8'h00;
14'h319e:data=8'h00;
14'h319f:data=8'h00;
14'h31a0:data=8'h1E;
14'h31a1:data=8'h00;
14'h31a2:data=8'h00;
14'h31a3:data=8'h00;
14'h31a4:data=8'h00;
14'h31a5:data=8'h00;
14'h31a6:data=8'h00;
14'h31a7:data=8'h00;
14'h31c0:data=8'h00;
14'h31c1:data=8'h00;
14'h31c2:data=8'h00;
14'h31c3:data=8'h00;
14'h31c4:data=8'h00;
14'h31c5:data=8'h00;
14'h31c6:data=8'h00;
14'h31c7:data=8'h00;
14'h31c8:data=8'h00;
14'h31c9:data=8'h07;
14'h31ca:data=8'hE0;
14'h31cb:data=8'h00;
14'h31cc:data=8'h00;
14'h31cd:data=8'h00;
14'h31ce:data=8'h00;
14'h31cf:data=8'h00;
14'h31d0:data=8'h00;
14'h31d1:data=8'h00;
14'h31d2:data=8'h03;
14'h31d3:data=8'hE0;
14'h31d4:data=8'h00;
14'h31d5:data=8'h00;
14'h31d6:data=8'h00;
14'h31d7:data=8'h00;
14'h31d8:data=8'h00;
14'h31d9:data=8'h00;
14'h31da:data=8'h00;
14'h31db:data=8'h00;
14'h31dc:data=8'h00;
14'h31dd:data=8'h00;
14'h31de:data=8'h00;
14'h31df:data=8'h03;
14'h31e0:data=8'hFC;
14'h31e1:data=8'h00;
14'h31e2:data=8'h00;
14'h31e3:data=8'h00;
14'h31e4:data=8'h00;
14'h31e5:data=8'h00;
14'h31e6:data=8'h00;
14'h31e7:data=8'h00;
14'h3200:data=8'h00;
14'h3201:data=8'h00;
14'h3202:data=8'h00;
14'h3203:data=8'h00;
14'h3204:data=8'h00;
14'h3205:data=8'h00;
14'h3206:data=8'h00;
14'h3207:data=8'h00;
14'h3208:data=8'h00;
14'h3209:data=8'hF8;
14'h320a:data=8'h00;
14'h320b:data=8'h00;
14'h320c:data=8'h00;
14'h320d:data=8'h00;
14'h320e:data=8'h00;
14'h320f:data=8'h00;
14'h3210:data=8'h00;
14'h3211:data=8'h00;
14'h3212:data=8'h7C;
14'h3213:data=8'h00;
14'h3214:data=8'h00;
14'h3215:data=8'h00;
14'h3216:data=8'h00;
14'h3217:data=8'h00;
14'h3218:data=8'h00;
14'h3219:data=8'h00;
14'h321a:data=8'h00;
14'h321b:data=8'h00;
14'h321c:data=8'h00;
14'h321d:data=8'h00;
14'h321e:data=8'h00;
14'h321f:data=8'h3F;
14'h3220:data=8'hFE;
14'h3221:data=8'h00;
14'h3222:data=8'h00;
14'h3223:data=8'h00;
14'h3224:data=8'h00;
14'h3225:data=8'h00;
14'h3226:data=8'h00;
14'h3227:data=8'h00;
14'h3240:data=8'h00;
14'h3241:data=8'h00;
14'h3242:data=8'h00;
14'h3243:data=8'h00;
14'h3244:data=8'h00;
14'h3245:data=8'h00;
14'h3246:data=8'h00;
14'h3247:data=8'h00;
14'h3248:data=8'h1F;
14'h3249:data=8'h00;
14'h324a:data=8'h00;
14'h324b:data=8'h00;
14'h324c:data=8'h00;
14'h324d:data=8'h00;
14'h324e:data=8'h00;
14'h324f:data=8'h00;
14'h3250:data=8'h00;
14'h3251:data=8'h0F;
14'h3252:data=8'h80;
14'h3253:data=8'h00;
14'h3254:data=8'h00;
14'h3255:data=8'h00;
14'h3256:data=8'h00;
14'h3257:data=8'h00;
14'h3258:data=8'h00;
14'h3259:data=8'h00;
14'h325a:data=8'h00;
14'h325b:data=8'h00;
14'h325c:data=8'h00;
14'h325d:data=8'h00;
14'h325e:data=8'h03;
14'h325f:data=8'hFF;
14'h3260:data=8'hFE;
14'h3261:data=8'h00;
14'h3262:data=8'h00;
14'h3263:data=8'h00;
14'h3264:data=8'h00;
14'h3265:data=8'h00;
14'h3266:data=8'h00;
14'h3267:data=8'h00;
14'h3280:data=8'h00;
14'h3281:data=8'h00;
14'h3282:data=8'h00;
14'h3283:data=8'h00;
14'h3284:data=8'h00;
14'h3285:data=8'h00;
14'h3286:data=8'h00;
14'h3287:data=8'h03;
14'h3288:data=8'hE0;
14'h3289:data=8'h00;
14'h328a:data=8'h00;
14'h328b:data=8'h00;
14'h328c:data=8'h00;
14'h328d:data=8'h00;
14'h328e:data=8'h00;
14'h328f:data=8'h00;
14'h3290:data=8'h01;
14'h3291:data=8'hF0;
14'h3292:data=8'h00;
14'h3293:data=8'h00;
14'h3294:data=8'h00;
14'h3295:data=8'h00;
14'h3296:data=8'h00;
14'h3297:data=8'h00;
14'h3298:data=8'h00;
14'h3299:data=8'h00;
14'h329a:data=8'h00;
14'h329b:data=8'h00;
14'h329c:data=8'h00;
14'h329d:data=8'h00;
14'h329e:data=8'h7F;
14'h329f:data=8'hFF;
14'h32a0:data=8'hFE;
14'h32a1:data=8'h00;
14'h32a2:data=8'h00;
14'h32a3:data=8'h00;
14'h32a4:data=8'h00;
14'h32a5:data=8'h00;
14'h32a6:data=8'h00;
14'h32a7:data=8'h00;
14'h32c0:data=8'h00;
14'h32c1:data=8'h00;
14'h32c2:data=8'h00;
14'h32c3:data=8'h00;
14'h32c4:data=8'h00;
14'h32c5:data=8'h00;
14'h32c6:data=8'h01;
14'h32c7:data=8'hFE;
14'h32c8:data=8'h00;
14'h32c9:data=8'h00;
14'h32ca:data=8'h00;
14'h32cb:data=8'h00;
14'h32cc:data=8'h00;
14'h32cd:data=8'h00;
14'h32ce:data=8'h00;
14'h32cf:data=8'h00;
14'h32d0:data=8'h3E;
14'h32d1:data=8'h00;
14'h32d2:data=8'h00;
14'h32d3:data=8'h00;
14'h32d4:data=8'h00;
14'h32d5:data=8'h00;
14'h32d6:data=8'h00;
14'h32d7:data=8'h00;
14'h32d8:data=8'h00;
14'h32d9:data=8'h00;
14'h32da:data=8'h00;
14'h32db:data=8'h00;
14'h32dc:data=8'h00;
14'h32dd:data=8'h07;
14'h32de:data=8'hFF;
14'h32df:data=8'hFF;
14'h32e0:data=8'hFE;
14'h32e1:data=8'h00;
14'h32e2:data=8'h00;
14'h32e3:data=8'h00;
14'h32e4:data=8'h00;
14'h32e5:data=8'h00;
14'h32e6:data=8'h00;
14'h32e7:data=8'h00;
14'h3300:data=8'h00;
14'h3301:data=8'h00;
14'h3302:data=8'h00;
14'h3303:data=8'h00;
14'h3304:data=8'h1F;
14'h3305:data=8'hFF;
14'h3306:data=8'hFF;
14'h3307:data=8'h00;
14'h3308:data=8'h00;
14'h3309:data=8'h00;
14'h330a:data=8'h00;
14'h330b:data=8'h00;
14'h330c:data=8'h00;
14'h330d:data=8'h00;
14'h330e:data=8'h00;
14'h330f:data=8'h0F;
14'h3310:data=8'hC0;
14'h3311:data=8'h00;
14'h3312:data=8'h00;
14'h3313:data=8'h00;
14'h3314:data=8'h00;
14'h3315:data=8'h00;
14'h3316:data=8'h00;
14'h3317:data=8'h00;
14'h3318:data=8'h00;
14'h3319:data=8'h00;
14'h331a:data=8'h00;
14'h331b:data=8'h00;
14'h331c:data=8'h00;
14'h331d:data=8'hFF;
14'h331e:data=8'hFF;
14'h331f:data=8'hFF;
14'h3320:data=8'hFE;
14'h3321:data=8'h00;
14'h3322:data=8'h00;
14'h3323:data=8'h00;
14'h3324:data=8'h00;
14'h3325:data=8'h00;
14'h3326:data=8'h00;
14'h3327:data=8'h00;
14'h3340:data=8'h00;
14'h3341:data=8'h00;
14'h3342:data=8'hFF;
14'h3343:data=8'hFF;
14'h3344:data=8'hF8;
14'h3345:data=8'h00;
14'h3346:data=8'h00;
14'h3347:data=8'h00;
14'h3348:data=8'h00;
14'h3349:data=8'h00;
14'h334a:data=8'h00;
14'h334b:data=8'h00;
14'h334c:data=8'h00;
14'h334d:data=8'h00;
14'h334e:data=8'h01;
14'h334f:data=8'hF8;
14'h3350:data=8'h00;
14'h3351:data=8'h00;
14'h3352:data=8'h00;
14'h3353:data=8'h00;
14'h3354:data=8'h00;
14'h3355:data=8'h00;
14'h3356:data=8'h00;
14'h3357:data=8'h00;
14'h3358:data=8'h00;
14'h3359:data=8'h00;
14'h335a:data=8'h00;
14'h335b:data=8'h00;
14'h335c:data=8'h0F;
14'h335d:data=8'hFF;
14'h335e:data=8'hFF;
14'h335f:data=8'hFF;
14'h3360:data=8'hFE;
14'h3361:data=8'h00;
14'h3362:data=8'h00;
14'h3363:data=8'h00;
14'h3364:data=8'h00;
14'h3365:data=8'h00;
14'h3366:data=8'h00;
14'h3367:data=8'h00;
14'h3380:data=8'hFF;
14'h3381:data=8'hFF;
14'h3382:data=8'h80;
14'h3383:data=8'h00;
14'h3384:data=8'h00;
14'h3385:data=8'h00;
14'h3386:data=8'h00;
14'h3387:data=8'h00;
14'h3388:data=8'h00;
14'h3389:data=8'h00;
14'h338a:data=8'h00;
14'h338b:data=8'h00;
14'h338c:data=8'h00;
14'h338d:data=8'h00;
14'h338e:data=8'h1F;
14'h338f:data=8'h00;
14'h3390:data=8'h00;
14'h3391:data=8'h00;
14'h3392:data=8'h00;
14'h3393:data=8'h00;
14'h3394:data=8'h00;
14'h3395:data=8'h00;
14'h3396:data=8'h00;
14'h3397:data=8'h00;
14'h3398:data=8'h00;
14'h3399:data=8'h00;
14'h339a:data=8'h00;
14'h339b:data=8'h00;
14'h339c:data=8'hFF;
14'h339d:data=8'hFF;
14'h339e:data=8'hFF;
14'h339f:data=8'hFF;
14'h33a0:data=8'hFE;
14'h33a1:data=8'h00;
14'h33a2:data=8'h00;
14'h33a3:data=8'h00;
14'h33a4:data=8'h00;
14'h33a5:data=8'h00;
14'h33a6:data=8'h00;
14'h33a7:data=8'h00;
14'h33c0:data=8'h00;
14'h33c1:data=8'h00;
14'h33c2:data=8'h00;
14'h33c3:data=8'h00;
14'h33c4:data=8'h00;
14'h33c5:data=8'h00;
14'h33c6:data=8'h00;
14'h33c7:data=8'h00;
14'h33c8:data=8'h00;
14'h33c9:data=8'h00;
14'h33ca:data=8'h00;
14'h33cb:data=8'h00;
14'h33cc:data=8'h00;
14'h33cd:data=8'h03;
14'h33ce:data=8'hE0;
14'h33cf:data=8'h00;
14'h33d0:data=8'h00;
14'h33d1:data=8'h00;
14'h33d2:data=8'h00;
14'h33d3:data=8'h00;
14'h33d4:data=8'h00;
14'h33d5:data=8'h00;
14'h33d6:data=8'h00;
14'h33d7:data=8'h00;
14'h33d8:data=8'h00;
14'h33d9:data=8'h00;
14'h33da:data=8'h00;
14'h33db:data=8'h0F;
14'h33dc:data=8'hFF;
14'h33dd:data=8'hFF;
14'h33de:data=8'hFF;
14'h33df:data=8'hFF;
14'h33e0:data=8'hFE;
14'h33e1:data=8'h00;
14'h33e2:data=8'h00;
14'h33e3:data=8'h00;
14'h33e4:data=8'h00;
14'h33e5:data=8'h00;
14'h33e6:data=8'h00;
14'h33e7:data=8'h00;
14'h3400:data=8'h00;
14'h3401:data=8'h00;
14'h3402:data=8'h00;
14'h3403:data=8'h00;
14'h3404:data=8'h00;
14'h3405:data=8'h00;
14'h3406:data=8'h00;
14'h3407:data=8'h00;
14'h3408:data=8'h00;
14'h3409:data=8'h00;
14'h340a:data=8'h00;
14'h340b:data=8'h00;
14'h340c:data=8'h00;
14'h340d:data=8'hF0;
14'h340e:data=8'h00;
14'h340f:data=8'h00;
14'h3410:data=8'h00;
14'h3411:data=8'h00;
14'h3412:data=8'h00;
14'h3413:data=8'h00;
14'h3414:data=8'h00;
14'h3415:data=8'h00;
14'h3416:data=8'h00;
14'h3417:data=8'h00;
14'h3418:data=8'h00;
14'h3419:data=8'h00;
14'h341a:data=8'h01;
14'h341b:data=8'hFF;
14'h341c:data=8'hFF;
14'h341d:data=8'hFF;
14'h341e:data=8'hFF;
14'h341f:data=8'hFF;
14'h3420:data=8'hFE;
14'h3421:data=8'h00;
14'h3422:data=8'h00;
14'h3423:data=8'h00;
14'h3424:data=8'h00;
14'h3425:data=8'h00;
14'h3426:data=8'h00;
14'h3427:data=8'h00;
14'h3440:data=8'h00;
14'h3441:data=8'h00;
14'h3442:data=8'h00;
14'h3443:data=8'h00;
14'h3444:data=8'h00;
14'h3445:data=8'h00;
14'h3446:data=8'h00;
14'h3447:data=8'h00;
14'h3448:data=8'h00;
14'h3449:data=8'h00;
14'h344a:data=8'h00;
14'h344b:data=8'h00;
14'h344c:data=8'h1E;
14'h344d:data=8'h00;
14'h344e:data=8'h00;
14'h344f:data=8'h00;
14'h3450:data=8'h00;
14'h3451:data=8'h00;
14'h3452:data=8'h00;
14'h3453:data=8'h00;
14'h3454:data=8'h00;
14'h3455:data=8'h00;
14'h3456:data=8'h00;
14'h3457:data=8'h00;
14'h3458:data=8'h00;
14'h3459:data=8'h00;
14'h345a:data=8'h01;
14'h345b:data=8'hFF;
14'h345c:data=8'hFF;
14'h345d:data=8'hFF;
14'h345e:data=8'hFF;
14'h345f:data=8'hFF;
14'h3460:data=8'hFE;
14'h3461:data=8'h00;
14'h3462:data=8'h00;
14'h3463:data=8'h00;
14'h3464:data=8'h00;
14'h3465:data=8'h00;
14'h3466:data=8'h00;
14'h3467:data=8'h00;
14'h3480:data=8'h00;
14'h3481:data=8'h00;
14'h3482:data=8'h00;
14'h3483:data=8'h00;
14'h3484:data=8'h00;
14'h3485:data=8'h00;
14'h3486:data=8'h00;
14'h3487:data=8'h00;
14'h3488:data=8'h00;
14'h3489:data=8'h00;
14'h348a:data=8'h00;
14'h348b:data=8'h03;
14'h348c:data=8'hC0;
14'h348d:data=8'h00;
14'h348e:data=8'h00;
14'h348f:data=8'h00;
14'h3490:data=8'h00;
14'h3491:data=8'h00;
14'h3492:data=8'h00;
14'h3493:data=8'h00;
14'h3494:data=8'h00;
14'h3495:data=8'h00;
14'h3496:data=8'h00;
14'h3497:data=8'h00;
14'h3498:data=8'h00;
14'h3499:data=8'h00;
14'h349a:data=8'h01;
14'h349b:data=8'hFF;
14'h349c:data=8'hFF;
14'h349d:data=8'hFF;
14'h349e:data=8'hFF;
14'h349f:data=8'hFF;
14'h34a0:data=8'hFE;
14'h34a1:data=8'h00;
14'h34a2:data=8'h00;
14'h34a3:data=8'h00;
14'h34a4:data=8'h00;
14'h34a5:data=8'h00;
14'h34a6:data=8'h00;
14'h34a7:data=8'h00;
14'h34c0:data=8'h00;
14'h34c1:data=8'h00;
14'h34c2:data=8'h00;
14'h34c3:data=8'h00;
14'h34c4:data=8'h00;
14'h34c5:data=8'h00;
14'h34c6:data=8'h00;
14'h34c7:data=8'h00;
14'h34c8:data=8'h00;
14'h34c9:data=8'h00;
14'h34ca:data=8'h00;
14'h34cb:data=8'h78;
14'h34cc:data=8'h00;
14'h34cd:data=8'h00;
14'h34ce:data=8'h00;
14'h34cf:data=8'h00;
14'h34d0:data=8'h00;
14'h34d1:data=8'h00;
14'h34d2:data=8'h00;
14'h34d3:data=8'h00;
14'h34d4:data=8'h00;
14'h34d5:data=8'h00;
14'h34d6:data=8'h00;
14'h34d7:data=8'h00;
14'h34d8:data=8'h00;
14'h34d9:data=8'h00;
14'h34da:data=8'h01;
14'h34db:data=8'hFF;
14'h34dc:data=8'hFF;
14'h34dd:data=8'hFF;
14'h34de:data=8'hFF;
14'h34df:data=8'hFF;
14'h34e0:data=8'hFE;
14'h34e1:data=8'h00;
14'h34e2:data=8'h00;
14'h34e3:data=8'h7F;
14'h34e4:data=8'hF0;
14'h34e5:data=8'h00;
14'h34e6:data=8'h00;
14'h34e7:data=8'h00;
14'h3500:data=8'h00;
14'h3501:data=8'h00;
14'h3502:data=8'h00;
14'h3503:data=8'h00;
14'h3504:data=8'h00;
14'h3505:data=8'h00;
14'h3506:data=8'h00;
14'h3507:data=8'h00;
14'h3508:data=8'h00;
14'h3509:data=8'h00;
14'h350a:data=8'h1F;
14'h350b:data=8'h00;
14'h350c:data=8'h00;
14'h350d:data=8'h00;
14'h350e:data=8'h00;
14'h350f:data=8'h00;
14'h3510:data=8'h00;
14'h3511:data=8'h00;
14'h3512:data=8'h00;
14'h3513:data=8'h00;
14'h3514:data=8'h00;
14'h3515:data=8'h00;
14'h3516:data=8'h00;
14'h3517:data=8'h00;
14'h3518:data=8'h00;
14'h3519:data=8'h00;
14'h351a:data=8'h01;
14'h351b:data=8'hFF;
14'h351c:data=8'hFF;
14'h351d:data=8'hFF;
14'h351e:data=8'hFF;
14'h351f:data=8'hFF;
14'h3520:data=8'hFE;
14'h3521:data=8'h00;
14'h3522:data=8'h00;
14'h3523:data=8'h7F;
14'h3524:data=8'hF0;
14'h3525:data=8'h00;
14'h3526:data=8'h00;
14'h3527:data=8'h00;
14'h3540:data=8'h00;
14'h3541:data=8'h00;
14'h3542:data=8'h00;
14'h3543:data=8'h00;
14'h3544:data=8'h00;
14'h3545:data=8'h00;
14'h3546:data=8'h00;
14'h3547:data=8'h00;
14'h3548:data=8'h00;
14'h3549:data=8'h03;
14'h354a:data=8'hC0;
14'h354b:data=8'h00;
14'h354c:data=8'h00;
14'h354d:data=8'h00;
14'h354e:data=8'h00;
14'h354f:data=8'h00;
14'h3550:data=8'h00;
14'h3551:data=8'h00;
14'h3552:data=8'h00;
14'h3553:data=8'h00;
14'h3554:data=8'h00;
14'h3555:data=8'h00;
14'h3556:data=8'h00;
14'h3557:data=8'h00;
14'h3558:data=8'h00;
14'h3559:data=8'h00;
14'h355a:data=8'h01;
14'h355b:data=8'hFF;
14'h355c:data=8'hFF;
14'h355d:data=8'hFF;
14'h355e:data=8'hFF;
14'h355f:data=8'hFF;
14'h3560:data=8'hFE;
14'h3561:data=8'h00;
14'h3562:data=8'h00;
14'h3563:data=8'h7F;
14'h3564:data=8'hF0;
14'h3565:data=8'h00;
14'h3566:data=8'h00;
14'h3567:data=8'h00;
14'h3580:data=8'h00;
14'h3581:data=8'h00;
14'h3582:data=8'h00;
14'h3583:data=8'h00;
14'h3584:data=8'h00;
14'h3585:data=8'h00;
14'h3586:data=8'h00;
14'h3587:data=8'h00;
14'h3588:data=8'h00;
14'h3589:data=8'h78;
14'h358a:data=8'h00;
14'h358b:data=8'h00;
14'h358c:data=8'h00;
14'h358d:data=8'h00;
14'h358e:data=8'h00;
14'h358f:data=8'h00;
14'h3590:data=8'h00;
14'h3591:data=8'h00;
14'h3592:data=8'h00;
14'h3593:data=8'h00;
14'h3594:data=8'h00;
14'h3595:data=8'h00;
14'h3596:data=8'h00;
14'h3597:data=8'h00;
14'h3598:data=8'h00;
14'h3599:data=8'h00;
14'h359a:data=8'h01;
14'h359b:data=8'hFF;
14'h359c:data=8'hFF;
14'h359d:data=8'hFF;
14'h359e:data=8'hFF;
14'h359f:data=8'hFF;
14'h35a0:data=8'hFF;
14'h35a1:data=8'h00;
14'h35a2:data=8'h00;
14'h35a3:data=8'h7F;
14'h35a4:data=8'hFF;
14'h35a5:data=8'hFE;
14'h35a6:data=8'h00;
14'h35a7:data=8'h00;
14'h35c0:data=8'h00;
14'h35c1:data=8'h00;
14'h35c2:data=8'h00;
14'h35c3:data=8'h00;
14'h35c4:data=8'h00;
14'h35c5:data=8'h00;
14'h35c6:data=8'h00;
14'h35c7:data=8'h00;
14'h35c8:data=8'h0F;
14'h35c9:data=8'h00;
14'h35ca:data=8'h00;
14'h35cb:data=8'h00;
14'h35cc:data=8'h00;
14'h35cd:data=8'h00;
14'h35ce:data=8'h00;
14'h35cf:data=8'h00;
14'h35d0:data=8'h00;
14'h35d1:data=8'h00;
14'h35d2:data=8'h00;
14'h35d3:data=8'h00;
14'h35d4:data=8'h00;
14'h35d5:data=8'h00;
14'h35d6:data=8'h00;
14'h35d7:data=8'h00;
14'h35d8:data=8'h00;
14'h35d9:data=8'h00;
14'h35da:data=8'h01;
14'h35db:data=8'hFF;
14'h35dc:data=8'hFF;
14'h35dd:data=8'hFF;
14'h35de:data=8'hFF;
14'h35df:data=8'hFF;
14'h35e0:data=8'hFF;
14'h35e1:data=8'h00;
14'h35e2:data=8'h00;
14'h35e3:data=8'h7F;
14'h35e4:data=8'hFF;
14'h35e5:data=8'hFE;
14'h35e6:data=8'h00;
14'h35e7:data=8'h00;
14'h3600:data=8'h00;
14'h3601:data=8'h00;
14'h3602:data=8'h00;
14'h3603:data=8'h00;
14'h3604:data=8'h00;
14'h3605:data=8'h00;
14'h3606:data=8'h00;
14'h3607:data=8'h07;
14'h3608:data=8'hE0;
14'h3609:data=8'h00;
14'h360a:data=8'h00;
14'h360b:data=8'h00;
14'h360c:data=8'h00;
14'h360d:data=8'h00;
14'h360e:data=8'h00;
14'h360f:data=8'h00;
14'h3610:data=8'h00;
14'h3611:data=8'h00;
14'h3612:data=8'h00;
14'h3613:data=8'h00;
14'h3614:data=8'h00;
14'h3615:data=8'h00;
14'h3616:data=8'h00;
14'h3617:data=8'h00;
14'h3618:data=8'h00;
14'h3619:data=8'h00;
14'h361a:data=8'h01;
14'h361b:data=8'hFF;
14'h361c:data=8'hFF;
14'h361d:data=8'hFF;
14'h361e:data=8'hFF;
14'h361f:data=8'hFF;
14'h3620:data=8'hFF;
14'h3621:data=8'h00;
14'h3622:data=8'h00;
14'h3623:data=8'h7F;
14'h3624:data=8'hFF;
14'h3625:data=8'hFE;
14'h3626:data=8'h00;
14'h3627:data=8'h00;
14'h3640:data=8'h00;
14'h3641:data=8'h00;
14'h3642:data=8'h00;
14'h3643:data=8'h00;
14'h3644:data=8'h03;
14'h3645:data=8'hFF;
14'h3646:data=8'hFF;
14'h3647:data=8'h80;
14'h3648:data=8'h00;
14'h3649:data=8'h00;
14'h364a:data=8'h00;
14'h364b:data=8'h00;
14'h364c:data=8'h00;
14'h364d:data=8'h00;
14'h364e:data=8'h00;
14'h364f:data=8'h00;
14'h3650:data=8'h00;
14'h3651:data=8'h00;
14'h3652:data=8'h00;
14'h3653:data=8'h00;
14'h3654:data=8'h00;
14'h3655:data=8'h00;
14'h3656:data=8'h00;
14'h3657:data=8'h00;
14'h3658:data=8'h00;
14'h3659:data=8'h00;
14'h365a:data=8'h01;
14'h365b:data=8'hFF;
14'h365c:data=8'hFF;
14'h365d:data=8'hFF;
14'h365e:data=8'hFF;
14'h365f:data=8'hFF;
14'h3660:data=8'hFF;
14'h3661:data=8'h00;
14'h3662:data=8'h00;
14'h3663:data=8'h7F;
14'h3664:data=8'hFF;
14'h3665:data=8'hFE;
14'h3666:data=8'h00;
14'h3667:data=8'h00;
14'h3680:data=8'h00;
14'h3681:data=8'h00;
14'h3682:data=8'h07;
14'h3683:data=8'hFF;
14'h3684:data=8'hFE;
14'h3685:data=8'h00;
14'h3686:data=8'h00;
14'h3687:data=8'h00;
14'h3688:data=8'h00;
14'h3689:data=8'h00;
14'h368a:data=8'h00;
14'h368b:data=8'h00;
14'h368c:data=8'h00;
14'h368d:data=8'h00;
14'h368e:data=8'h00;
14'h368f:data=8'h00;
14'h3690:data=8'h00;
14'h3691:data=8'h00;
14'h3692:data=8'h00;
14'h3693:data=8'h00;
14'h3694:data=8'h00;
14'h3695:data=8'h00;
14'h3696:data=8'h00;
14'h3697:data=8'h00;
14'h3698:data=8'h00;
14'h3699:data=8'h00;
14'h369a:data=8'h01;
14'h369b:data=8'hFF;
14'h369c:data=8'hFF;
14'h369d:data=8'hFF;
14'h369e:data=8'hFF;
14'h369f:data=8'hFF;
14'h36a0:data=8'hFF;
14'h36a1:data=8'h00;
14'h36a2:data=8'h00;
14'h36a3:data=8'h7F;
14'h36a4:data=8'hFF;
14'h36a5:data=8'hFE;
14'h36a6:data=8'h00;
14'h36a7:data=8'h00;
14'h36c0:data=8'h1F;
14'h36c1:data=8'hFF;
14'h36c2:data=8'hFC;
14'h36c3:data=8'h00;
14'h36c4:data=8'h00;
14'h36c5:data=8'h00;
14'h36c6:data=8'h00;
14'h36c7:data=8'h00;
14'h36c8:data=8'h00;
14'h36c9:data=8'h00;
14'h36ca:data=8'h00;
14'h36cb:data=8'h00;
14'h36cc:data=8'h00;
14'h36cd:data=8'h00;
14'h36ce:data=8'h00;
14'h36cf:data=8'h00;
14'h36d0:data=8'h00;
14'h36d1:data=8'h00;
14'h36d2:data=8'h00;
14'h36d3:data=8'h00;
14'h36d4:data=8'h00;
14'h36d5:data=8'h00;
14'h36d6:data=8'h00;
14'h36d7:data=8'h00;
14'h36d8:data=8'h00;
14'h36d9:data=8'h00;
14'h36da:data=8'h01;
14'h36db:data=8'hFF;
14'h36dc:data=8'hFF;
14'h36dd:data=8'hFF;
14'h36de:data=8'hFF;
14'h36df:data=8'hFF;
14'h36e0:data=8'hFF;
14'h36e1:data=8'h00;
14'h36e2:data=8'h00;
14'h36e3:data=8'h7F;
14'h36e4:data=8'hFF;
14'h36e5:data=8'hFE;
14'h36e6:data=8'h00;
14'h36e7:data=8'h00;
14'h3700:data=8'hF0;
14'h3701:data=8'h00;
14'h3702:data=8'h00;
14'h3703:data=8'h00;
14'h3704:data=8'h00;
14'h3705:data=8'h00;
14'h3706:data=8'h00;
14'h3707:data=8'h00;
14'h3708:data=8'h00;
14'h3709:data=8'h00;
14'h370a:data=8'h00;
14'h370b:data=8'h00;
14'h370c:data=8'h00;
14'h370d:data=8'h00;
14'h370e:data=8'h00;
14'h370f:data=8'h00;
14'h3710:data=8'h00;
14'h3711:data=8'h00;
14'h3712:data=8'h00;
14'h3713:data=8'h00;
14'h3714:data=8'h00;
14'h3715:data=8'h00;
14'h3716:data=8'h00;
14'h3717:data=8'h00;
14'h3718:data=8'h00;
14'h3719:data=8'h00;
14'h371a:data=8'h01;
14'h371b:data=8'hFF;
14'h371c:data=8'hFF;
14'h371d:data=8'hFF;
14'h371e:data=8'hFF;
14'h371f:data=8'hFF;
14'h3720:data=8'hFF;
14'h3721:data=8'hFF;
14'h3722:data=8'hFF;
14'h3723:data=8'hFF;
14'h3724:data=8'hFF;
14'h3725:data=8'hFE;
14'h3726:data=8'h00;
14'h3727:data=8'h00;
14'h3740:data=8'h00;
14'h3741:data=8'h00;
14'h3742:data=8'h00;
14'h3743:data=8'h00;
14'h3744:data=8'h00;
14'h3745:data=8'h00;
14'h3746:data=8'h00;
14'h3747:data=8'h00;
14'h3748:data=8'h00;
14'h3749:data=8'h00;
14'h374a:data=8'h00;
14'h374b:data=8'h00;
14'h374c:data=8'h00;
14'h374d:data=8'h00;
14'h374e:data=8'h00;
14'h374f:data=8'h00;
14'h3750:data=8'h00;
14'h3751:data=8'h00;
14'h3752:data=8'h00;
14'h3753:data=8'h00;
14'h3754:data=8'h00;
14'h3755:data=8'h00;
14'h3756:data=8'h00;
14'h3757:data=8'h00;
14'h3758:data=8'h00;
14'h3759:data=8'h00;
14'h375a:data=8'h01;
14'h375b:data=8'hFF;
14'h375c:data=8'hFF;
14'h375d:data=8'hFF;
14'h375e:data=8'hFF;
14'h375f:data=8'hFF;
14'h3760:data=8'hFF;
14'h3761:data=8'hFF;
14'h3762:data=8'hFF;
14'h3763:data=8'hFF;
14'h3764:data=8'hFF;
14'h3765:data=8'hFE;
14'h3766:data=8'h00;
14'h3767:data=8'h00;
14'h3780:data=8'h00;
14'h3781:data=8'h00;
14'h3782:data=8'h00;
14'h3783:data=8'h00;
14'h3784:data=8'h00;
14'h3785:data=8'h00;
14'h3786:data=8'h00;
14'h3787:data=8'h00;
14'h3788:data=8'h00;
14'h3789:data=8'h00;
14'h378a:data=8'h00;
14'h378b:data=8'h00;
14'h378c:data=8'h00;
14'h378d:data=8'h00;
14'h378e:data=8'h00;
14'h378f:data=8'h00;
14'h3790:data=8'h00;
14'h3791:data=8'h00;
14'h3792:data=8'h00;
14'h3793:data=8'h00;
14'h3794:data=8'h00;
14'h3795:data=8'h00;
14'h3796:data=8'h00;
14'h3797:data=8'h00;
14'h3798:data=8'h00;
14'h3799:data=8'h00;
14'h379a:data=8'h01;
14'h379b:data=8'hFF;
14'h379c:data=8'hFF;
14'h379d:data=8'hFF;
14'h379e:data=8'hFF;
14'h379f:data=8'hFF;
14'h37a0:data=8'hFF;
14'h37a1:data=8'hFF;
14'h37a2:data=8'hFF;
14'h37a3:data=8'hFF;
14'h37a4:data=8'hFF;
14'h37a5:data=8'hFE;
14'h37a6:data=8'h00;
14'h37a7:data=8'h00;
14'h37c0:data=8'h00;
14'h37c1:data=8'h00;
14'h37c2:data=8'h00;
14'h37c3:data=8'h00;
14'h37c4:data=8'h00;
14'h37c5:data=8'h00;
14'h37c6:data=8'h00;
14'h37c7:data=8'h00;
14'h37c8:data=8'h00;
14'h37c9:data=8'h00;
14'h37ca:data=8'h00;
14'h37cb:data=8'h00;
14'h37cc:data=8'h00;
14'h37cd:data=8'h00;
14'h37ce:data=8'h00;
14'h37cf:data=8'h00;
14'h37d0:data=8'h00;
14'h37d1:data=8'h00;
14'h37d2:data=8'h00;
14'h37d3:data=8'h00;
14'h37d4:data=8'h00;
14'h37d5:data=8'h00;
14'h37d6:data=8'h00;
14'h37d7:data=8'h00;
14'h37d8:data=8'h00;
14'h37d9:data=8'h00;
14'h37da:data=8'h01;
14'h37db:data=8'hFF;
14'h37dc:data=8'hFF;
14'h37dd:data=8'hFF;
14'h37de:data=8'hFF;
14'h37df:data=8'hFF;
14'h37e0:data=8'hFF;
14'h37e1:data=8'hFF;
14'h37e2:data=8'hFF;
14'h37e3:data=8'hFF;
14'h37e4:data=8'hFF;
14'h37e5:data=8'hFE;
14'h37e6:data=8'h00;
14'h37e7:data=8'h00;
14'h3800:data=8'h00;
14'h3801:data=8'h00;
14'h3802:data=8'h00;
14'h3803:data=8'h00;
14'h3804:data=8'h00;
14'h3805:data=8'h00;
14'h3806:data=8'h00;
14'h3807:data=8'h00;
14'h3808:data=8'h00;
14'h3809:data=8'h00;
14'h380a:data=8'h00;
14'h380b:data=8'h00;
14'h380c:data=8'h00;
14'h380d:data=8'h00;
14'h380e:data=8'h00;
14'h380f:data=8'h00;
14'h3810:data=8'h00;
14'h3811:data=8'h00;
14'h3812:data=8'h00;
14'h3813:data=8'h00;
14'h3814:data=8'h00;
14'h3815:data=8'h00;
14'h3816:data=8'h00;
14'h3817:data=8'h00;
14'h3818:data=8'h00;
14'h3819:data=8'h00;
14'h381a:data=8'h01;
14'h381b:data=8'hFF;
14'h381c:data=8'hFF;
14'h381d:data=8'hFF;
14'h381e:data=8'hFF;
14'h381f:data=8'hFF;
14'h3820:data=8'hFF;
14'h3821:data=8'hFF;
14'h3822:data=8'hFF;
14'h3823:data=8'hFF;
14'h3824:data=8'hFF;
14'h3825:data=8'hFF;
14'h3826:data=8'h00;
14'h3827:data=8'h00;
14'h3840:data=8'h00;
14'h3841:data=8'h00;
14'h3842:data=8'h00;
14'h3843:data=8'h00;
14'h3844:data=8'h00;
14'h3845:data=8'h00;
14'h3846:data=8'h00;
14'h3847:data=8'h00;
14'h3848:data=8'h00;
14'h3849:data=8'h00;
14'h384a:data=8'h00;
14'h384b:data=8'h00;
14'h384c:data=8'h00;
14'h384d:data=8'h00;
14'h384e:data=8'h00;
14'h384f:data=8'h00;
14'h3850:data=8'h00;
14'h3851:data=8'h00;
14'h3852:data=8'h00;
14'h3853:data=8'h00;
14'h3854:data=8'h00;
14'h3855:data=8'h00;
14'h3856:data=8'h00;
14'h3857:data=8'h00;
14'h3858:data=8'h00;
14'h3859:data=8'h00;
14'h385a:data=8'h01;
14'h385b:data=8'hFF;
14'h385c:data=8'hFF;
14'h385d:data=8'hFF;
14'h385e:data=8'hFF;
14'h385f:data=8'hFF;
14'h3860:data=8'hFF;
14'h3861:data=8'hFF;
14'h3862:data=8'hFF;
14'h3863:data=8'hFF;
14'h3864:data=8'hFF;
14'h3865:data=8'hFF;
14'h3866:data=8'h00;
14'h3867:data=8'h00;
14'h3880:data=8'h00;
14'h3881:data=8'h00;
14'h3882:data=8'h00;
14'h3883:data=8'h00;
14'h3884:data=8'h00;
14'h3885:data=8'h00;
14'h3886:data=8'h00;
14'h3887:data=8'h00;
14'h3888:data=8'h00;
14'h3889:data=8'h00;
14'h388a:data=8'h00;
14'h388b:data=8'h00;
14'h388c:data=8'h00;
14'h388d:data=8'h00;
14'h388e:data=8'h00;
14'h388f:data=8'h00;
14'h3890:data=8'h00;
14'h3891:data=8'h00;
14'h3892:data=8'h00;
14'h3893:data=8'h00;
14'h3894:data=8'h00;
14'h3895:data=8'h00;
14'h3896:data=8'h00;
14'h3897:data=8'h00;
14'h3898:data=8'h00;
14'h3899:data=8'h00;
14'h389a:data=8'h01;
14'h389b:data=8'hFF;
14'h389c:data=8'hFF;
14'h389d:data=8'hFF;
14'h389e:data=8'hFF;
14'h389f:data=8'hFF;
14'h38a0:data=8'hFF;
14'h38a1:data=8'hFF;
14'h38a2:data=8'hFF;
14'h38a3:data=8'hFF;
14'h38a4:data=8'hFF;
14'h38a5:data=8'hFF;
14'h38a6:data=8'h00;
14'h38a7:data=8'h00;
14'h38c0:data=8'h00;
14'h38c1:data=8'h00;
14'h38c2:data=8'h00;
14'h38c3:data=8'h00;
14'h38c4:data=8'h00;
14'h38c5:data=8'h00;
14'h38c6:data=8'h00;
14'h38c7:data=8'h00;
14'h38c8:data=8'h00;
14'h38c9:data=8'h00;
14'h38ca:data=8'h00;
14'h38cb:data=8'h00;
14'h38cc:data=8'h00;
14'h38cd:data=8'h00;
14'h38ce:data=8'h00;
14'h38cf:data=8'h00;
14'h38d0:data=8'h00;
14'h38d1:data=8'h00;
14'h38d2:data=8'h00;
14'h38d3:data=8'h00;
14'h38d4:data=8'h00;
14'h38d5:data=8'h00;
14'h38d6:data=8'h00;
14'h38d7:data=8'h00;
14'h38d8:data=8'h00;
14'h38d9:data=8'h00;
14'h38da:data=8'h01;
14'h38db:data=8'hFF;
14'h38dc:data=8'hFF;
14'h38dd:data=8'hFF;
14'h38de:data=8'hFF;
14'h38df:data=8'hFF;
14'h38e0:data=8'hFF;
14'h38e1:data=8'hFF;
14'h38e2:data=8'hFF;
14'h38e3:data=8'hFF;
14'h38e4:data=8'hFF;
14'h38e5:data=8'hFF;
14'h38e6:data=8'h00;
14'h38e7:data=8'h00;
14'h3900:data=8'h00;
14'h3901:data=8'h00;
14'h3902:data=8'h00;
14'h3903:data=8'h00;
14'h3904:data=8'h00;
14'h3905:data=8'h00;
14'h3906:data=8'h00;
14'h3907:data=8'h00;
14'h3908:data=8'h00;
14'h3909:data=8'h00;
14'h390a:data=8'h00;
14'h390b:data=8'h00;
14'h390c:data=8'h00;
14'h390d:data=8'h00;
14'h390e:data=8'h00;
14'h390f:data=8'h00;
14'h3910:data=8'h00;
14'h3911:data=8'h00;
14'h3912:data=8'h00;
14'h3913:data=8'h00;
14'h3914:data=8'h00;
14'h3915:data=8'h00;
14'h3916:data=8'h00;
14'h3917:data=8'h00;
14'h3918:data=8'h00;
14'h3919:data=8'h00;
14'h391a:data=8'h01;
14'h391b:data=8'hFF;
14'h391c:data=8'hFF;
14'h391d:data=8'hFF;
14'h391e:data=8'hFF;
14'h391f:data=8'hFF;
14'h3920:data=8'hFF;
14'h3921:data=8'hFF;
14'h3922:data=8'hFF;
14'h3923:data=8'hFF;
14'h3924:data=8'hFF;
14'h3925:data=8'hFF;
14'h3926:data=8'h00;
14'h3927:data=8'h00;
14'h3940:data=8'h00;
14'h3941:data=8'h00;
14'h3942:data=8'h00;
14'h3943:data=8'h00;
14'h3944:data=8'h00;
14'h3945:data=8'h00;
14'h3946:data=8'h00;
14'h3947:data=8'h00;
14'h3948:data=8'h00;
14'h3949:data=8'h00;
14'h394a:data=8'h00;
14'h394b:data=8'h00;
14'h394c:data=8'h00;
14'h394d:data=8'h00;
14'h394e:data=8'h00;
14'h394f:data=8'h00;
14'h3950:data=8'h00;
14'h3951:data=8'h00;
14'h3952:data=8'h00;
14'h3953:data=8'h00;
14'h3954:data=8'h00;
14'h3955:data=8'h00;
14'h3956:data=8'h00;
14'h3957:data=8'h00;
14'h3958:data=8'h00;
14'h3959:data=8'h00;
14'h395a:data=8'h01;
14'h395b:data=8'hFF;
14'h395c:data=8'hFF;
14'h395d:data=8'hFF;
14'h395e:data=8'hFF;
14'h395f:data=8'hFE;
14'h3960:data=8'h00;
14'h3961:data=8'h00;
14'h3962:data=8'h00;
14'h3963:data=8'h3F;
14'h3964:data=8'hFF;
14'h3965:data=8'hFF;
14'h3966:data=8'h00;
14'h3967:data=8'h00;
14'h3980:data=8'h00;
14'h3981:data=8'h00;
14'h3982:data=8'h00;
14'h3983:data=8'h00;
14'h3984:data=8'h00;
14'h3985:data=8'h00;
14'h3986:data=8'h00;
14'h3987:data=8'h00;
14'h3988:data=8'h00;
14'h3989:data=8'h00;
14'h398a:data=8'h00;
14'h398b:data=8'h00;
14'h398c:data=8'h00;
14'h398d:data=8'h00;
14'h398e:data=8'h00;
14'h398f:data=8'h00;
14'h3990:data=8'h00;
14'h3991:data=8'h00;
14'h3992:data=8'h00;
14'h3993:data=8'h00;
14'h3994:data=8'h00;
14'h3995:data=8'h00;
14'h3996:data=8'h00;
14'h3997:data=8'h00;
14'h3998:data=8'h00;
14'h3999:data=8'h00;
14'h399a:data=8'h01;
14'h399b:data=8'hFF;
14'h399c:data=8'hFF;
14'h399d:data=8'hFF;
14'h399e:data=8'hFF;
14'h399f:data=8'hFE;
14'h39a0:data=8'h00;
14'h39a1:data=8'h00;
14'h39a2:data=8'h00;
14'h39a3:data=8'h3F;
14'h39a4:data=8'hFF;
14'h39a5:data=8'hFF;
14'h39a6:data=8'h00;
14'h39a7:data=8'h00;
14'h39c0:data=8'h00;
14'h39c1:data=8'h00;
14'h39c2:data=8'h00;
14'h39c3:data=8'h00;
14'h39c4:data=8'h00;
14'h39c5:data=8'h00;
14'h39c6:data=8'h00;
14'h39c7:data=8'h00;
14'h39c8:data=8'h00;
14'h39c9:data=8'h00;
14'h39ca:data=8'h00;
14'h39cb:data=8'h00;
14'h39cc:data=8'h00;
14'h39cd:data=8'h00;
14'h39ce:data=8'h00;
14'h39cf:data=8'h00;
14'h39d0:data=8'h00;
14'h39d1:data=8'h00;
14'h39d2:data=8'h00;
14'h39d3:data=8'h00;
14'h39d4:data=8'h00;
14'h39d5:data=8'h00;
14'h39d6:data=8'h00;
14'h39d7:data=8'h00;
14'h39d8:data=8'h00;
14'h39d9:data=8'h00;
14'h39da:data=8'h01;
14'h39db:data=8'hFF;
14'h39dc:data=8'hFF;
14'h39dd:data=8'hFF;
14'h39de:data=8'hFF;
14'h39df:data=8'hFE;
14'h39e0:data=8'h00;
14'h39e1:data=8'h00;
14'h39e2:data=8'h00;
14'h39e3:data=8'h3F;
14'h39e4:data=8'hFF;
14'h39e5:data=8'hFF;
14'h39e6:data=8'h00;
14'h39e7:data=8'h00;
14'h3a00:data=8'h00;
14'h3a01:data=8'h00;
14'h3a02:data=8'h00;
14'h3a03:data=8'h00;
14'h3a04:data=8'h00;
14'h3a05:data=8'h00;
14'h3a06:data=8'h00;
14'h3a07:data=8'h00;
14'h3a08:data=8'h00;
14'h3a09:data=8'h00;
14'h3a0a:data=8'h00;
14'h3a0b:data=8'h00;
14'h3a0c:data=8'h00;
14'h3a0d:data=8'h00;
14'h3a0e:data=8'h00;
14'h3a0f:data=8'h00;
14'h3a10:data=8'h00;
14'h3a11:data=8'h00;
14'h3a12:data=8'h00;
14'h3a13:data=8'h00;
14'h3a14:data=8'h00;
14'h3a15:data=8'h00;
14'h3a16:data=8'h00;
14'h3a17:data=8'h00;
14'h3a18:data=8'h00;
14'h3a19:data=8'h00;
14'h3a1a:data=8'h01;
14'h3a1b:data=8'hFF;
14'h3a1c:data=8'hFF;
14'h3a1d:data=8'hFF;
14'h3a1e:data=8'hFF;
14'h3a1f:data=8'hFE;
14'h3a20:data=8'h00;
14'h3a21:data=8'h00;
14'h3a22:data=8'h00;
14'h3a23:data=8'h3F;
14'h3a24:data=8'hFF;
14'h3a25:data=8'hFF;
14'h3a26:data=8'h00;
14'h3a27:data=8'h00;
14'h3a40:data=8'h00;
14'h3a41:data=8'h00;
14'h3a42:data=8'h00;
14'h3a43:data=8'h00;
14'h3a44:data=8'h00;
14'h3a45:data=8'h00;
14'h3a46:data=8'h00;
14'h3a47:data=8'h00;
14'h3a48:data=8'h00;
14'h3a49:data=8'h00;
14'h3a4a:data=8'h00;
14'h3a4b:data=8'h00;
14'h3a4c:data=8'h00;
14'h3a4d:data=8'h00;
14'h3a4e:data=8'h00;
14'h3a4f:data=8'h00;
14'h3a50:data=8'h00;
14'h3a51:data=8'h00;
14'h3a52:data=8'h00;
14'h3a53:data=8'h00;
14'h3a54:data=8'h00;
14'h3a55:data=8'h00;
14'h3a56:data=8'h00;
14'h3a57:data=8'h00;
14'h3a58:data=8'h00;
14'h3a59:data=8'h00;
14'h3a5a:data=8'h01;
14'h3a5b:data=8'hFF;
14'h3a5c:data=8'hFF;
14'h3a5d:data=8'hFF;
14'h3a5e:data=8'hFF;
14'h3a5f:data=8'hFE;
14'h3a60:data=8'h00;
14'h3a61:data=8'h00;
14'h3a62:data=8'h00;
14'h3a63:data=8'h3F;
14'h3a64:data=8'hFF;
14'h3a65:data=8'hFF;
14'h3a66:data=8'h00;
14'h3a67:data=8'h00;
14'h3a80:data=8'h00;
14'h3a81:data=8'h00;
14'h3a82:data=8'h00;
14'h3a83:data=8'h00;
14'h3a84:data=8'h00;
14'h3a85:data=8'h00;
14'h3a86:data=8'h00;
14'h3a87:data=8'h00;
14'h3a88:data=8'h00;
14'h3a89:data=8'h00;
14'h3a8a:data=8'h00;
14'h3a8b:data=8'h00;
14'h3a8c:data=8'h00;
14'h3a8d:data=8'h00;
14'h3a8e:data=8'h00;
14'h3a8f:data=8'h00;
14'h3a90:data=8'h00;
14'h3a91:data=8'h00;
14'h3a92:data=8'h00;
14'h3a93:data=8'h00;
14'h3a94:data=8'h00;
14'h3a95:data=8'h00;
14'h3a96:data=8'h00;
14'h3a97:data=8'h00;
14'h3a98:data=8'h00;
14'h3a99:data=8'h00;
14'h3a9a:data=8'h01;
14'h3a9b:data=8'hFF;
14'h3a9c:data=8'hFF;
14'h3a9d:data=8'hFF;
14'h3a9e:data=8'hFF;
14'h3a9f:data=8'hFE;
14'h3aa0:data=8'h00;
14'h3aa1:data=8'h00;
14'h3aa2:data=8'h00;
14'h3aa3:data=8'h3F;
14'h3aa4:data=8'hFF;
14'h3aa5:data=8'hFF;
14'h3aa6:data=8'h00;
14'h3aa7:data=8'h00;
14'h3ac0:data=8'h00;
14'h3ac1:data=8'h00;
14'h3ac2:data=8'h00;
14'h3ac3:data=8'h00;
14'h3ac4:data=8'h00;
14'h3ac5:data=8'h00;
14'h3ac6:data=8'h00;
14'h3ac7:data=8'h00;
14'h3ac8:data=8'h00;
14'h3ac9:data=8'h00;
14'h3aca:data=8'h00;
14'h3acb:data=8'h00;
14'h3acc:data=8'h00;
14'h3acd:data=8'h00;
14'h3ace:data=8'h00;
14'h3acf:data=8'h00;
14'h3ad0:data=8'h00;
14'h3ad1:data=8'h00;
14'h3ad2:data=8'h00;
14'h3ad3:data=8'h00;
14'h3ad4:data=8'h00;
14'h3ad5:data=8'h00;
14'h3ad6:data=8'h00;
14'h3ad7:data=8'h00;
14'h3ad8:data=8'h00;
14'h3ad9:data=8'h00;
14'h3ada:data=8'h01;
14'h3adb:data=8'hFF;
14'h3adc:data=8'hFF;
14'h3add:data=8'hFF;
14'h3ade:data=8'hFF;
14'h3adf:data=8'hFE;
14'h3ae0:data=8'h00;
14'h3ae1:data=8'h00;
14'h3ae2:data=8'h00;
14'h3ae3:data=8'h3F;
14'h3ae4:data=8'hFF;
14'h3ae5:data=8'hFF;
14'h3ae6:data=8'h00;
14'h3ae7:data=8'h00;
14'h3b00:data=8'h00;
14'h3b01:data=8'h00;
14'h3b02:data=8'h00;
14'h3b03:data=8'h00;
14'h3b04:data=8'h00;
14'h3b05:data=8'h00;
14'h3b06:data=8'h00;
14'h3b07:data=8'h00;
14'h3b08:data=8'h00;
14'h3b09:data=8'h00;
14'h3b0a:data=8'h00;
14'h3b0b:data=8'h00;
14'h3b0c:data=8'h00;
14'h3b0d:data=8'h00;
14'h3b0e:data=8'h00;
14'h3b0f:data=8'h00;
14'h3b10:data=8'h00;
14'h3b11:data=8'h00;
14'h3b12:data=8'h00;
14'h3b13:data=8'h00;
14'h3b14:data=8'h00;
14'h3b15:data=8'h00;
14'h3b16:data=8'h00;
14'h3b17:data=8'h00;
14'h3b18:data=8'h00;
14'h3b19:data=8'h00;
14'h3b1a:data=8'h01;
14'h3b1b:data=8'hFF;
14'h3b1c:data=8'hFF;
14'h3b1d:data=8'hFF;
14'h3b1e:data=8'hFF;
14'h3b1f:data=8'hFE;
14'h3b20:data=8'h00;
14'h3b21:data=8'h00;
14'h3b22:data=8'h00;
14'h3b23:data=8'h3F;
14'h3b24:data=8'hFF;
14'h3b25:data=8'hFF;
14'h3b26:data=8'h00;
14'h3b27:data=8'h00;
14'h3b40:data=8'h00;
14'h3b41:data=8'h00;
14'h3b42:data=8'h00;
14'h3b43:data=8'h00;
14'h3b44:data=8'h00;
14'h3b45:data=8'h00;
14'h3b46:data=8'h00;
14'h3b47:data=8'h00;
14'h3b48:data=8'h00;
14'h3b49:data=8'h00;
14'h3b4a:data=8'h00;
14'h3b4b:data=8'h00;
14'h3b4c:data=8'h00;
14'h3b4d:data=8'h00;
14'h3b4e:data=8'h00;
14'h3b4f:data=8'h00;
14'h3b50:data=8'h00;
14'h3b51:data=8'h00;
14'h3b52:data=8'h00;
14'h3b53:data=8'h00;
14'h3b54:data=8'h00;
14'h3b55:data=8'h00;
14'h3b56:data=8'h00;
14'h3b57:data=8'h00;
14'h3b58:data=8'h00;
14'h3b59:data=8'h00;
14'h3b5a:data=8'h01;
14'h3b5b:data=8'hFF;
14'h3b5c:data=8'hFF;
14'h3b5d:data=8'hFF;
14'h3b5e:data=8'hFF;
14'h3b5f:data=8'hFE;
14'h3b60:data=8'h00;
14'h3b61:data=8'h00;
14'h3b62:data=8'h00;
14'h3b63:data=8'h3F;
14'h3b64:data=8'hFF;
14'h3b65:data=8'hFF;
14'h3b66:data=8'h00;
14'h3b67:data=8'h00;
14'h3b80:data=8'h00;
14'h3b81:data=8'h00;
14'h3b82:data=8'h00;
14'h3b83:data=8'h00;
14'h3b84:data=8'h00;
14'h3b85:data=8'h00;
14'h3b86:data=8'h00;
14'h3b87:data=8'h00;
14'h3b88:data=8'h00;
14'h3b89:data=8'h00;
14'h3b8a:data=8'h00;
14'h3b8b:data=8'h00;
14'h3b8c:data=8'h00;
14'h3b8d:data=8'h00;
14'h3b8e:data=8'h00;
14'h3b8f:data=8'h00;
14'h3b90:data=8'h00;
14'h3b91:data=8'h00;
14'h3b92:data=8'h00;
14'h3b93:data=8'h00;
14'h3b94:data=8'h00;
14'h3b95:data=8'h00;
14'h3b96:data=8'h00;
14'h3b97:data=8'h00;
14'h3b98:data=8'h00;
14'h3b99:data=8'h00;
14'h3b9a:data=8'h01;
14'h3b9b:data=8'hFF;
14'h3b9c:data=8'hFF;
14'h3b9d:data=8'hFF;
14'h3b9e:data=8'hFF;
14'h3b9f:data=8'hFE;
14'h3ba0:data=8'h00;
14'h3ba1:data=8'h00;
14'h3ba2:data=8'h00;
14'h3ba3:data=8'h3F;
14'h3ba4:data=8'hFF;
14'h3ba5:data=8'hFF;
14'h3ba6:data=8'h00;
14'h3ba7:data=8'h00;
14'h3bc0:data=8'hff;
14'h3bc1:data=8'hff;
14'h3bc2:data=8'hff;
14'h3bc3:data=8'hff;
14'h3bc4:data=8'hff;
14'h3bc5:data=8'hff;
14'h3bc6:data=8'hff;
14'h3bc7:data=8'hff;
14'h3bc8:data=8'hff;
14'h3bc9:data=8'hff;
14'h3bca:data=8'hff;
14'h3bcb:data=8'hff;
14'h3bcc:data=8'hff;
14'h3bcd:data=8'hff;
14'h3bce:data=8'hff;
14'h3bcf:data=8'hff;
14'h3bd0:data=8'hff;
14'h3bd1:data=8'hff;
14'h3bd2:data=8'hff;
14'h3bd3:data=8'hff;
14'h3bd4:data=8'hff;
14'h3bd5:data=8'hff;
14'h3bd6:data=8'hff;
14'h3bd7:data=8'hff;
14'h3bd8:data=8'hff;
14'h3bd9:data=8'hff;
14'h3bda:data=8'hff;
14'h3bdb:data=8'hff;
14'h3bdc:data=8'hff;
14'h3bdd:data=8'hff;
14'h3bde:data=8'hff;
14'h3bdf:data=8'hff;
14'h3be0:data=8'hff;
14'h3be1:data=8'hff;
14'h3be2:data=8'hff;
14'h3be3:data=8'hff;
14'h3be4:data=8'hff;
14'h3be5:data=8'hff;
14'h3be6:data=8'hff;
14'h3be7:data=8'hff;

			
		default:data=8'h00;
		endcase
	end
endmodule
