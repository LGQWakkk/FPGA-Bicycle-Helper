`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/06/15 16:16:31
// Design Name: 
// Module Name: big_digit_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//20230615 19:16 V1
//20230615 20:31 V1 测试成功（改正了显示顺序反的问题）
module big_digit_rom(
	input wire clk,
	input wire [14:0] addr,//15bit addr
	output reg [7:0] data
    );
	
	//数据结构：{[6:0],[2:0],[4:0]} {ASCII[6:0],ROW[2:0],COL_24[4:0]}
	//ASCII:0X30-0X39  ROW:0-5!!!!!  COL:0-23
	reg [14:0] addr_reg;
	
	always@(posedge clk)begin
		addr_reg<=addr;
	end
	
	always@(*)begin
		case(addr_reg)
15'h3000:data=8'h00;
15'h3001:data=8'h00;
15'h3002:data=8'h00;
15'h3003:data=8'h00;
15'h3004:data=8'h00;
15'h3005:data=8'h00;
15'h3006:data=8'h00;
15'h3007:data=8'h00;
15'h3008:data=8'h00;
15'h3009:data=8'h00;
15'h300a:data=8'h00;
15'h300b:data=8'h80;
15'h300c:data=8'h80;
15'h300d:data=8'h00;
15'h300e:data=8'h00;
15'h300f:data=8'h00;
15'h3010:data=8'h00;
15'h3011:data=8'h00;
15'h3012:data=8'h00;
15'h3013:data=8'h00;
15'h3014:data=8'h00;
15'h3015:data=8'h00;
15'h3016:data=8'h00;
15'h3017:data=8'h00;
15'h3020:data=8'h00;
15'h3021:data=8'h00;
15'h3022:data=8'h00;
15'h3023:data=8'hE0;
15'h3024:data=8'hF0;
15'h3025:data=8'hFC;
15'h3026:data=8'hFE;
15'h3027:data=8'h3E;
15'h3028:data=8'h1F;
15'h3029:data=8'h0F;
15'h302a:data=8'h07;
15'h302b:data=8'h07;
15'h302c:data=8'h07;
15'h302d:data=8'h07;
15'h302e:data=8'h0F;
15'h302f:data=8'h1F;
15'h3030:data=8'h7E;
15'h3031:data=8'hFC;
15'h3032:data=8'hF8;
15'h3033:data=8'hE0;
15'h3034:data=8'h80;
15'h3035:data=8'h00;
15'h3036:data=8'h00;
15'h3037:data=8'h00;
15'h3040:data=8'h00;
15'h3041:data=8'h00;
15'h3042:data=8'hFF;
15'h3043:data=8'hFF;
15'h3044:data=8'hFF;
15'h3045:data=8'h3F;
15'h3046:data=8'h00;
15'h3047:data=8'h00;
15'h3048:data=8'h00;
15'h3049:data=8'h00;
15'h304a:data=8'h00;
15'h304b:data=8'h00;
15'h304c:data=8'h00;
15'h304d:data=8'h00;
15'h304e:data=8'h00;
15'h304f:data=8'h00;
15'h3050:data=8'h00;
15'h3051:data=8'h07;
15'h3052:data=8'hFF;
15'h3053:data=8'hFF;
15'h3054:data=8'hFF;
15'h3055:data=8'hC0;
15'h3056:data=8'h00;
15'h3057:data=8'h00;
15'h3060:data=8'h00;
15'h3061:data=8'h00;
15'h3062:data=8'hFF;
15'h3063:data=8'hFF;
15'h3064:data=8'hFF;
15'h3065:data=8'hF8;
15'h3066:data=8'h00;
15'h3067:data=8'h00;
15'h3068:data=8'h00;
15'h3069:data=8'h00;
15'h306a:data=8'h00;
15'h306b:data=8'h00;
15'h306c:data=8'h00;
15'h306d:data=8'h00;
15'h306e:data=8'h00;
15'h306f:data=8'h00;
15'h3070:data=8'h00;
15'h3071:data=8'hE0;
15'h3072:data=8'hFF;
15'h3073:data=8'hFF;
15'h3074:data=8'hFF;
15'h3075:data=8'h03;
15'h3076:data=8'h00;
15'h3077:data=8'h00;
15'h3080:data=8'h00;
15'h3081:data=8'h00;
15'h3082:data=8'h00;
15'h3083:data=8'h03;
15'h3084:data=8'h0F;
15'h3085:data=8'h3F;
15'h3086:data=8'h3F;
15'h3087:data=8'h7C;
15'h3088:data=8'hF8;
15'h3089:data=8'hF0;
15'h308a:data=8'hE0;
15'h308b:data=8'hE0;
15'h308c:data=8'hE0;
15'h308d:data=8'hF0;
15'h308e:data=8'hF0;
15'h308f:data=8'hF8;
15'h3090:data=8'h7E;
15'h3091:data=8'h3F;
15'h3092:data=8'h1F;
15'h3093:data=8'h07;
15'h3094:data=8'h01;
15'h3095:data=8'h00;
15'h3096:data=8'h00;
15'h3097:data=8'h00;
15'h30a0:data=8'h00;
15'h30a1:data=8'h00;
15'h30a2:data=8'h00;
15'h30a3:data=8'h00;
15'h30a4:data=8'h00;
15'h30a5:data=8'h00;
15'h30a6:data=8'h00;
15'h30a7:data=8'h00;
15'h30a8:data=8'h00;
15'h30a9:data=8'h00;
15'h30aa:data=8'h00;
15'h30ab:data=8'h00;
15'h30ac:data=8'h00;
15'h30ad:data=8'h00;
15'h30ae:data=8'h00;
15'h30af:data=8'h00;
15'h30b0:data=8'h00;
15'h30b1:data=8'h00;
15'h30b2:data=8'h00;
15'h30b3:data=8'h00;
15'h30b4:data=8'h00;
15'h30b5:data=8'h00;
15'h30b6:data=8'h00;
15'h30b7:data=8'h00;

15'h3100:data=8'h00;
15'h3101:data=8'h00;
15'h3102:data=8'h00;
15'h3103:data=8'h00;
15'h3104:data=8'h00;
15'h3105:data=8'h00;
15'h3106:data=8'h00;
15'h3107:data=8'h00;
15'h3108:data=8'h00;
15'h3109:data=8'h00;
15'h310a:data=8'h00;
15'h310b:data=8'h00;
15'h310c:data=8'h00;
15'h310d:data=8'h00;
15'h310e:data=8'h00;
15'h310f:data=8'h00;
15'h3110:data=8'h00;
15'h3111:data=8'h00;
15'h3112:data=8'h00;
15'h3113:data=8'h00;
15'h3114:data=8'h00;
15'h3115:data=8'h00;
15'h3116:data=8'h00;
15'h3117:data=8'h00;
15'h3120:data=8'h00;
15'h3121:data=8'h00;
15'h3122:data=8'h00;
15'h3123:data=8'h00;
15'h3124:data=8'h80;
15'h3125:data=8'hC0;
15'h3126:data=8'hC0;
15'h3127:data=8'hE0;
15'h3128:data=8'hF0;
15'h3129:data=8'h78;
15'h312a:data=8'hFC;
15'h312b:data=8'hFF;
15'h312c:data=8'hFF;
15'h312d:data=8'hFF;
15'h312e:data=8'h00;
15'h312f:data=8'h00;
15'h3130:data=8'h00;
15'h3131:data=8'h00;
15'h3132:data=8'h00;
15'h3133:data=8'h00;
15'h3134:data=8'h00;
15'h3135:data=8'h00;
15'h3136:data=8'h00;
15'h3137:data=8'h00;
15'h3140:data=8'h00;
15'h3141:data=8'h00;
15'h3142:data=8'h00;
15'h3143:data=8'h00;
15'h3144:data=8'h07;
15'h3145:data=8'h03;
15'h3146:data=8'h01;
15'h3147:data=8'h01;
15'h3148:data=8'h00;
15'h3149:data=8'h00;
15'h314a:data=8'hFF;
15'h314b:data=8'hFF;
15'h314c:data=8'hFF;
15'h314d:data=8'hFF;
15'h314e:data=8'h00;
15'h314f:data=8'h00;
15'h3150:data=8'h00;
15'h3151:data=8'h00;
15'h3152:data=8'h00;
15'h3153:data=8'h00;
15'h3154:data=8'h00;
15'h3155:data=8'h00;
15'h3156:data=8'h00;
15'h3157:data=8'h00;
15'h3160:data=8'h00;
15'h3161:data=8'h00;
15'h3162:data=8'h00;
15'h3163:data=8'h00;
15'h3164:data=8'h00;
15'h3165:data=8'h00;
15'h3166:data=8'h00;
15'h3167:data=8'h00;
15'h3168:data=8'h00;
15'h3169:data=8'h00;
15'h316a:data=8'hFF;
15'h316b:data=8'hFF;
15'h316c:data=8'hFF;
15'h316d:data=8'hFF;
15'h316e:data=8'h00;
15'h316f:data=8'h00;
15'h3170:data=8'h00;
15'h3171:data=8'h00;
15'h3172:data=8'h00;
15'h3173:data=8'h00;
15'h3174:data=8'h00;
15'h3175:data=8'h00;
15'h3176:data=8'h00;
15'h3177:data=8'h00;
15'h3180:data=8'h00;
15'h3181:data=8'h00;
15'h3182:data=8'h00;
15'h3183:data=8'h00;
15'h3184:data=8'h00;
15'h3185:data=8'h00;
15'h3186:data=8'h00;
15'h3187:data=8'h00;
15'h3188:data=8'h00;
15'h3189:data=8'h00;
15'h318a:data=8'hFF;
15'h318b:data=8'hFF;
15'h318c:data=8'hFF;
15'h318d:data=8'hFF;
15'h318e:data=8'h00;
15'h318f:data=8'h00;
15'h3190:data=8'h00;
15'h3191:data=8'h00;
15'h3192:data=8'h00;
15'h3193:data=8'h00;
15'h3194:data=8'h00;
15'h3195:data=8'h00;
15'h3196:data=8'h00;
15'h3197:data=8'h00;
15'h31a0:data=8'h00;
15'h31a1:data=8'h00;
15'h31a2:data=8'h00;
15'h31a3:data=8'h00;
15'h31a4:data=8'h00;
15'h31a5:data=8'h00;
15'h31a6:data=8'h00;
15'h31a7:data=8'h00;
15'h31a8:data=8'h00;
15'h31a9:data=8'h00;
15'h31aa:data=8'h00;
15'h31ab:data=8'h00;
15'h31ac:data=8'h00;
15'h31ad:data=8'h00;
15'h31ae:data=8'h00;
15'h31af:data=8'h00;
15'h31b0:data=8'h00;
15'h31b1:data=8'h00;
15'h31b2:data=8'h00;
15'h31b3:data=8'h00;
15'h31b4:data=8'h00;
15'h31b5:data=8'h00;
15'h31b6:data=8'h00;
15'h31b7:data=8'h00;

15'h3200:data=8'h00;
15'h3201:data=8'h00;
15'h3202:data=8'h00;
15'h3203:data=8'h00;
15'h3204:data=8'h00;
15'h3205:data=8'h00;
15'h3206:data=8'h00;
15'h3207:data=8'h00;
15'h3208:data=8'h00;
15'h3209:data=8'h00;
15'h320a:data=8'h80;
15'h320b:data=8'h80;
15'h320c:data=8'h80;
15'h320d:data=8'h80;
15'h320e:data=8'h00;
15'h320f:data=8'h00;
15'h3210:data=8'h00;
15'h3211:data=8'h00;
15'h3212:data=8'h00;
15'h3213:data=8'h00;
15'h3214:data=8'h00;
15'h3215:data=8'h00;
15'h3216:data=8'h00;
15'h3217:data=8'h00;
15'h3220:data=8'h00;
15'h3221:data=8'h00;
15'h3222:data=8'hE0;
15'h3223:data=8'hF0;
15'h3224:data=8'hFC;
15'h3225:data=8'h7E;
15'h3226:data=8'h3E;
15'h3227:data=8'h1F;
15'h3228:data=8'h0F;
15'h3229:data=8'h0F;
15'h322a:data=8'h07;
15'h322b:data=8'h07;
15'h322c:data=8'h07;
15'h322d:data=8'h07;
15'h322e:data=8'h0F;
15'h322f:data=8'h0F;
15'h3230:data=8'h3F;
15'h3231:data=8'hFE;
15'h3232:data=8'hFC;
15'h3233:data=8'hF8;
15'h3234:data=8'hE0;
15'h3235:data=8'h00;
15'h3236:data=8'h00;
15'h3237:data=8'h00;
15'h3240:data=8'h00;
15'h3241:data=8'h00;
15'h3242:data=8'h00;
15'h3243:data=8'h00;
15'h3244:data=8'h00;
15'h3245:data=8'h00;
15'h3246:data=8'h00;
15'h3247:data=8'h00;
15'h3248:data=8'h00;
15'h3249:data=8'h00;
15'h324a:data=8'h00;
15'h324b:data=8'h00;
15'h324c:data=8'h00;
15'h324d:data=8'h00;
15'h324e:data=8'hC0;
15'h324f:data=8'hE0;
15'h3250:data=8'hFC;
15'h3251:data=8'hFF;
15'h3252:data=8'h7F;
15'h3253:data=8'h1F;
15'h3254:data=8'h03;
15'h3255:data=8'h00;
15'h3256:data=8'h00;
15'h3257:data=8'h00;
15'h3260:data=8'h00;
15'h3261:data=8'h00;
15'h3262:data=8'h00;
15'h3263:data=8'h00;
15'h3264:data=8'h00;
15'h3265:data=8'h00;
15'h3266:data=8'h00;
15'h3267:data=8'h80;
15'h3268:data=8'hC0;
15'h3269:data=8'hE0;
15'h326a:data=8'hF0;
15'h326b:data=8'hFC;
15'h326c:data=8'h7E;
15'h326d:data=8'h3F;
15'h326e:data=8'h0F;
15'h326f:data=8'h07;
15'h3270:data=8'h03;
15'h3271:data=8'h00;
15'h3272:data=8'h00;
15'h3273:data=8'h00;
15'h3274:data=8'h00;
15'h3275:data=8'h00;
15'h3276:data=8'h00;
15'h3277:data=8'h00;
15'h3280:data=8'h00;
15'h3281:data=8'h00;
15'h3282:data=8'hC0;
15'h3283:data=8'hF0;
15'h3284:data=8'hFC;
15'h3285:data=8'hFE;
15'h3286:data=8'hFF;
15'h3287:data=8'hFF;
15'h3288:data=8'hFF;
15'h3289:data=8'hF3;
15'h328a:data=8'hF1;
15'h328b:data=8'hF0;
15'h328c:data=8'hF0;
15'h328d:data=8'hF0;
15'h328e:data=8'hF0;
15'h328f:data=8'hF0;
15'h3290:data=8'hF0;
15'h3291:data=8'hF0;
15'h3292:data=8'hF0;
15'h3293:data=8'hF0;
15'h3294:data=8'hF0;
15'h3295:data=8'h00;
15'h3296:data=8'h00;
15'h3297:data=8'h00;
15'h32a0:data=8'h00;
15'h32a1:data=8'h00;
15'h32a2:data=8'h00;
15'h32a3:data=8'h00;
15'h32a4:data=8'h00;
15'h32a5:data=8'h00;
15'h32a6:data=8'h00;
15'h32a7:data=8'h00;
15'h32a8:data=8'h00;
15'h32a9:data=8'h00;
15'h32aa:data=8'h00;
15'h32ab:data=8'h00;
15'h32ac:data=8'h00;
15'h32ad:data=8'h00;
15'h32ae:data=8'h00;
15'h32af:data=8'h00;
15'h32b0:data=8'h00;
15'h32b1:data=8'h00;
15'h32b2:data=8'h00;
15'h32b3:data=8'h00;
15'h32b4:data=8'h00;
15'h32b5:data=8'h00;
15'h32b6:data=8'h00;
15'h32b7:data=8'h00;

15'h3300:data=8'h00;
15'h3301:data=8'h00;
15'h3302:data=8'h00;
15'h3303:data=8'h00;
15'h3304:data=8'h00;
15'h3305:data=8'h00;
15'h3306:data=8'h00;
15'h3307:data=8'h00;
15'h3308:data=8'h00;
15'h3309:data=8'h00;
15'h330a:data=8'h00;
15'h330b:data=8'h00;
15'h330c:data=8'h00;
15'h330d:data=8'h00;
15'h330e:data=8'h00;
15'h330f:data=8'h00;
15'h3310:data=8'h00;
15'h3311:data=8'h00;
15'h3312:data=8'h00;
15'h3313:data=8'h00;
15'h3314:data=8'h00;
15'h3315:data=8'h00;
15'h3316:data=8'h00;
15'h3317:data=8'h00;
15'h3320:data=8'h00;
15'h3321:data=8'h00;
15'h3322:data=8'h80;
15'h3323:data=8'hE0;
15'h3324:data=8'hF8;
15'h3325:data=8'hFC;
15'h3326:data=8'h3E;
15'h3327:data=8'h1E;
15'h3328:data=8'h0F;
15'h3329:data=8'h07;
15'h332a:data=8'h07;
15'h332b:data=8'h07;
15'h332c:data=8'h07;
15'h332d:data=8'h07;
15'h332e:data=8'h0F;
15'h332f:data=8'h0F;
15'h3330:data=8'h3F;
15'h3331:data=8'hFE;
15'h3332:data=8'hFC;
15'h3333:data=8'hF8;
15'h3334:data=8'hE0;
15'h3335:data=8'h00;
15'h3336:data=8'h00;
15'h3337:data=8'h00;
15'h3340:data=8'h00;
15'h3341:data=8'h00;
15'h3342:data=8'h00;
15'h3343:data=8'h00;
15'h3344:data=8'h00;
15'h3345:data=8'h00;
15'h3346:data=8'h00;
15'h3347:data=8'h00;
15'h3348:data=8'h00;
15'h3349:data=8'h00;
15'h334a:data=8'hC0;
15'h334b:data=8'hC0;
15'h334c:data=8'hE0;
15'h334d:data=8'hE0;
15'h334e:data=8'hF0;
15'h334f:data=8'hF0;
15'h3350:data=8'hFC;
15'h3351:data=8'h3F;
15'h3352:data=8'h1F;
15'h3353:data=8'h0F;
15'h3354:data=8'h01;
15'h3355:data=8'h00;
15'h3356:data=8'h00;
15'h3357:data=8'h00;
15'h3360:data=8'h00;
15'h3361:data=8'h00;
15'h3362:data=8'h00;
15'h3363:data=8'h00;
15'h3364:data=8'h80;
15'h3365:data=8'h00;
15'h3366:data=8'h00;
15'h3367:data=8'h00;
15'h3368:data=8'h00;
15'h3369:data=8'h00;
15'h336a:data=8'h00;
15'h336b:data=8'h01;
15'h336c:data=8'h01;
15'h336d:data=8'h01;
15'h336e:data=8'h03;
15'h336f:data=8'h03;
15'h3370:data=8'h0F;
15'h3371:data=8'hFF;
15'h3372:data=8'hFF;
15'h3373:data=8'hFE;
15'h3374:data=8'hF8;
15'h3375:data=8'h00;
15'h3376:data=8'h00;
15'h3377:data=8'h00;
15'h3380:data=8'h00;
15'h3381:data=8'h00;
15'h3382:data=8'h03;
15'h3383:data=8'h0F;
15'h3384:data=8'h1F;
15'h3385:data=8'h3F;
15'h3386:data=8'h7C;
15'h3387:data=8'h78;
15'h3388:data=8'hF0;
15'h3389:data=8'hF0;
15'h338a:data=8'hE0;
15'h338b:data=8'hE0;
15'h338c:data=8'hE0;
15'h338d:data=8'hE0;
15'h338e:data=8'hF0;
15'h338f:data=8'hF8;
15'h3390:data=8'h7C;
15'h3391:data=8'h3F;
15'h3392:data=8'h3F;
15'h3393:data=8'h0F;
15'h3394:data=8'h07;
15'h3395:data=8'h00;
15'h3396:data=8'h00;
15'h3397:data=8'h00;
15'h33a0:data=8'h00;
15'h33a1:data=8'h00;
15'h33a2:data=8'h00;
15'h33a3:data=8'h00;
15'h33a4:data=8'h00;
15'h33a5:data=8'h00;
15'h33a6:data=8'h00;
15'h33a7:data=8'h00;
15'h33a8:data=8'h00;
15'h33a9:data=8'h00;
15'h33aa:data=8'h00;
15'h33ab:data=8'h00;
15'h33ac:data=8'h00;
15'h33ad:data=8'h00;
15'h33ae:data=8'h00;
15'h33af:data=8'h00;
15'h33b0:data=8'h00;
15'h33b1:data=8'h00;
15'h33b2:data=8'h00;
15'h33b3:data=8'h00;
15'h33b4:data=8'h00;
15'h33b5:data=8'h00;
15'h33b6:data=8'h00;
15'h33b7:data=8'h00;

15'h3400:data=8'h00;
15'h3401:data=8'h00;
15'h3402:data=8'h00;
15'h3403:data=8'h00;
15'h3404:data=8'h00;
15'h3405:data=8'h00;
15'h3406:data=8'h00;
15'h3407:data=8'h00;
15'h3408:data=8'h00;
15'h3409:data=8'h00;
15'h340a:data=8'h00;
15'h340b:data=8'h00;
15'h340c:data=8'h00;
15'h340d:data=8'h00;
15'h340e:data=8'h00;
15'h340f:data=8'h00;
15'h3410:data=8'h00;
15'h3411:data=8'h00;
15'h3412:data=8'h00;
15'h3413:data=8'h00;
15'h3414:data=8'h00;
15'h3415:data=8'h00;
15'h3416:data=8'h00;
15'h3417:data=8'h00;
15'h3420:data=8'h00;
15'h3421:data=8'h00;
15'h3422:data=8'h00;
15'h3423:data=8'h00;
15'h3424:data=8'h00;
15'h3425:data=8'h00;
15'h3426:data=8'h00;
15'h3427:data=8'h00;
15'h3428:data=8'h00;
15'h3429:data=8'h00;
15'h342a:data=8'h80;
15'h342b:data=8'hC0;
15'h342c:data=8'hF0;
15'h342d:data=8'hF8;
15'h342e:data=8'h7E;
15'h342f:data=8'hFF;
15'h3430:data=8'hFF;
15'h3431:data=8'hFF;
15'h3432:data=8'hFF;
15'h3433:data=8'h00;
15'h3434:data=8'h00;
15'h3435:data=8'h00;
15'h3436:data=8'h00;
15'h3437:data=8'h00;
15'h3440:data=8'h00;
15'h3441:data=8'h00;
15'h3442:data=8'h00;
15'h3443:data=8'h00;
15'h3444:data=8'h00;
15'h3445:data=8'hC0;
15'h3446:data=8'hE0;
15'h3447:data=8'hF0;
15'h3448:data=8'hFC;
15'h3449:data=8'h7E;
15'h344a:data=8'h1F;
15'h344b:data=8'h0F;
15'h344c:data=8'h03;
15'h344d:data=8'h01;
15'h344e:data=8'h00;
15'h344f:data=8'hFF;
15'h3450:data=8'hFF;
15'h3451:data=8'hFF;
15'h3452:data=8'hFF;
15'h3453:data=8'h00;
15'h3454:data=8'h00;
15'h3455:data=8'h00;
15'h3456:data=8'h00;
15'h3457:data=8'h00;
15'h3460:data=8'h00;
15'h3461:data=8'hF0;
15'h3462:data=8'hF8;
15'h3463:data=8'hFE;
15'h3464:data=8'hFF;
15'h3465:data=8'hCF;
15'h3466:data=8'hC7;
15'h3467:data=8'hC1;
15'h3468:data=8'hC0;
15'h3469:data=8'hC0;
15'h346a:data=8'hC0;
15'h346b:data=8'hC0;
15'h346c:data=8'hC0;
15'h346d:data=8'hC0;
15'h346e:data=8'hC0;
15'h346f:data=8'hFF;
15'h3470:data=8'hFF;
15'h3471:data=8'hFF;
15'h3472:data=8'hFF;
15'h3473:data=8'hC0;
15'h3474:data=8'hC0;
15'h3475:data=8'hC0;
15'h3476:data=8'hC0;
15'h3477:data=8'h00;
15'h3480:data=8'h00;
15'h3481:data=8'h01;
15'h3482:data=8'h01;
15'h3483:data=8'h01;
15'h3484:data=8'h01;
15'h3485:data=8'h01;
15'h3486:data=8'h01;
15'h3487:data=8'h01;
15'h3488:data=8'h01;
15'h3489:data=8'h01;
15'h348a:data=8'h01;
15'h348b:data=8'h01;
15'h348c:data=8'h01;
15'h348d:data=8'h01;
15'h348e:data=8'h01;
15'h348f:data=8'hFF;
15'h3490:data=8'hFF;
15'h3491:data=8'hFF;
15'h3492:data=8'hFF;
15'h3493:data=8'h01;
15'h3494:data=8'h01;
15'h3495:data=8'h01;
15'h3496:data=8'h01;
15'h3497:data=8'h00;
15'h34a0:data=8'h00;
15'h34a1:data=8'h00;
15'h34a2:data=8'h00;
15'h34a3:data=8'h00;
15'h34a4:data=8'h00;
15'h34a5:data=8'h00;
15'h34a6:data=8'h00;
15'h34a7:data=8'h00;
15'h34a8:data=8'h00;
15'h34a9:data=8'h00;
15'h34aa:data=8'h00;
15'h34ab:data=8'h00;
15'h34ac:data=8'h00;
15'h34ad:data=8'h00;
15'h34ae:data=8'h00;
15'h34af:data=8'h00;
15'h34b0:data=8'h00;
15'h34b1:data=8'h00;
15'h34b2:data=8'h00;
15'h34b3:data=8'h00;
15'h34b4:data=8'h00;
15'h34b5:data=8'h00;
15'h34b6:data=8'h00;
15'h34b7:data=8'h00;

15'h3500:data=8'h00;
15'h3501:data=8'h00;
15'h3502:data=8'h00;
15'h3503:data=8'h00;
15'h3504:data=8'h00;
15'h3505:data=8'h00;
15'h3506:data=8'h00;
15'h3507:data=8'h00;
15'h3508:data=8'h00;
15'h3509:data=8'h00;
15'h350a:data=8'h00;
15'h350b:data=8'h00;
15'h350c:data=8'h00;
15'h350d:data=8'h00;
15'h350e:data=8'h00;
15'h350f:data=8'h00;
15'h3510:data=8'h00;
15'h3511:data=8'h00;
15'h3512:data=8'h00;
15'h3513:data=8'h00;
15'h3514:data=8'h00;
15'h3515:data=8'h00;
15'h3516:data=8'h00;
15'h3517:data=8'h00;
15'h3520:data=8'h00;
15'h3521:data=8'h00;
15'h3522:data=8'h00;
15'h3523:data=8'h00;
15'h3524:data=8'hF0;
15'h3525:data=8'hFF;
15'h3526:data=8'hFF;
15'h3527:data=8'h3F;
15'h3528:data=8'h0F;
15'h3529:data=8'h0F;
15'h352a:data=8'h0F;
15'h352b:data=8'h0F;
15'h352c:data=8'h0F;
15'h352d:data=8'h0F;
15'h352e:data=8'h0F;
15'h352f:data=8'h0F;
15'h3530:data=8'h0F;
15'h3531:data=8'h0F;
15'h3532:data=8'h0F;
15'h3533:data=8'h0F;
15'h3534:data=8'h00;
15'h3535:data=8'h00;
15'h3536:data=8'h00;
15'h3537:data=8'h00;
15'h3540:data=8'h00;
15'h3541:data=8'h00;
15'h3542:data=8'hE0;
15'h3543:data=8'hFF;
15'h3544:data=8'hFF;
15'h3545:data=8'hFF;
15'h3546:data=8'h7F;
15'h3547:data=8'h38;
15'h3548:data=8'h38;
15'h3549:data=8'h38;
15'h354a:data=8'h3C;
15'h354b:data=8'h3C;
15'h354c:data=8'h3C;
15'h354d:data=8'h38;
15'h354e:data=8'h78;
15'h354f:data=8'hF8;
15'h3550:data=8'hF0;
15'h3551:data=8'hF0;
15'h3552:data=8'hE0;
15'h3553:data=8'h80;
15'h3554:data=8'h00;
15'h3555:data=8'h00;
15'h3556:data=8'h00;
15'h3557:data=8'h00;
15'h3560:data=8'h00;
15'h3561:data=8'h00;
15'h3562:data=8'h00;
15'h3563:data=8'h81;
15'h3564:data=8'h01;
15'h3565:data=8'h00;
15'h3566:data=8'h00;
15'h3567:data=8'h00;
15'h3568:data=8'h00;
15'h3569:data=8'h00;
15'h356a:data=8'h00;
15'h356b:data=8'h00;
15'h356c:data=8'h00;
15'h356d:data=8'h00;
15'h356e:data=8'h00;
15'h356f:data=8'h00;
15'h3570:data=8'h01;
15'h3571:data=8'hFF;
15'h3572:data=8'hFF;
15'h3573:data=8'hFF;
15'h3574:data=8'hFE;
15'h3575:data=8'h00;
15'h3576:data=8'h00;
15'h3577:data=8'h00;
15'h3580:data=8'h00;
15'h3581:data=8'h07;
15'h3582:data=8'h1F;
15'h3583:data=8'h3F;
15'h3584:data=8'h7F;
15'h3585:data=8'h7C;
15'h3586:data=8'hF0;
15'h3587:data=8'hF0;
15'h3588:data=8'hE0;
15'h3589:data=8'hE0;
15'h358a:data=8'hE0;
15'h358b:data=8'hE0;
15'h358c:data=8'hE0;
15'h358d:data=8'hF0;
15'h358e:data=8'hF0;
15'h358f:data=8'h78;
15'h3590:data=8'h7E;
15'h3591:data=8'h3F;
15'h3592:data=8'h1F;
15'h3593:data=8'h0F;
15'h3594:data=8'h03;
15'h3595:data=8'h00;
15'h3596:data=8'h00;
15'h3597:data=8'h00;
15'h35a0:data=8'h00;
15'h35a1:data=8'h00;
15'h35a2:data=8'h00;
15'h35a3:data=8'h00;
15'h35a4:data=8'h00;
15'h35a5:data=8'h00;
15'h35a6:data=8'h00;
15'h35a7:data=8'h00;
15'h35a8:data=8'h00;
15'h35a9:data=8'h00;
15'h35aa:data=8'h00;
15'h35ab:data=8'h00;
15'h35ac:data=8'h00;
15'h35ad:data=8'h00;
15'h35ae:data=8'h00;
15'h35af:data=8'h00;
15'h35b0:data=8'h00;
15'h35b1:data=8'h00;
15'h35b2:data=8'h00;
15'h35b3:data=8'h00;
15'h35b4:data=8'h00;
15'h35b5:data=8'h00;
15'h35b6:data=8'h00;
15'h35b7:data=8'h00;

15'h3600:data=8'h00;
15'h3601:data=8'h00;
15'h3602:data=8'h00;
15'h3603:data=8'h00;
15'h3604:data=8'h00;
15'h3605:data=8'h00;
15'h3606:data=8'h00;
15'h3607:data=8'h00;
15'h3608:data=8'h00;
15'h3609:data=8'h00;
15'h360a:data=8'h00;
15'h360b:data=8'h00;
15'h360c:data=8'h00;
15'h360d:data=8'h00;
15'h360e:data=8'h00;
15'h360f:data=8'h00;
15'h3610:data=8'h00;
15'h3611:data=8'h00;
15'h3612:data=8'h00;
15'h3613:data=8'h00;
15'h3614:data=8'h00;
15'h3615:data=8'h00;
15'h3616:data=8'h00;
15'h3617:data=8'h00;
15'h3620:data=8'h00;
15'h3621:data=8'h00;
15'h3622:data=8'h00;
15'h3623:data=8'h00;
15'h3624:data=8'h00;
15'h3625:data=8'h00;
15'h3626:data=8'h00;
15'h3627:data=8'h00;
15'h3628:data=8'h80;
15'h3629:data=8'hE0;
15'h362a:data=8'hF0;
15'h362b:data=8'hFC;
15'h362c:data=8'h7E;
15'h362d:data=8'h3F;
15'h362e:data=8'h0F;
15'h362f:data=8'h07;
15'h3630:data=8'h01;
15'h3631:data=8'h00;
15'h3632:data=8'h00;
15'h3633:data=8'h00;
15'h3634:data=8'h00;
15'h3635:data=8'h00;
15'h3636:data=8'h00;
15'h3637:data=8'h00;
15'h3640:data=8'h00;
15'h3641:data=8'h00;
15'h3642:data=8'h00;
15'h3643:data=8'h80;
15'h3644:data=8'hE0;
15'h3645:data=8'hF0;
15'h3646:data=8'hFC;
15'h3647:data=8'hFF;
15'h3648:data=8'hFF;
15'h3649:data=8'h7F;
15'h364a:data=8'h77;
15'h364b:data=8'h71;
15'h364c:data=8'h78;
15'h364d:data=8'h78;
15'h364e:data=8'h78;
15'h364f:data=8'h70;
15'h3650:data=8'hF0;
15'h3651:data=8'hF0;
15'h3652:data=8'hE0;
15'h3653:data=8'hC0;
15'h3654:data=8'h80;
15'h3655:data=8'h00;
15'h3656:data=8'h00;
15'h3657:data=8'h00;
15'h3660:data=8'h00;
15'h3661:data=8'h00;
15'h3662:data=8'hFE;
15'h3663:data=8'hFF;
15'h3664:data=8'hFF;
15'h3665:data=8'hFF;
15'h3666:data=8'h03;
15'h3667:data=8'h01;
15'h3668:data=8'h00;
15'h3669:data=8'h00;
15'h366a:data=8'h00;
15'h366b:data=8'h00;
15'h366c:data=8'h00;
15'h366d:data=8'h00;
15'h366e:data=8'h00;
15'h366f:data=8'h00;
15'h3670:data=8'h00;
15'h3671:data=8'h01;
15'h3672:data=8'h07;
15'h3673:data=8'hFF;
15'h3674:data=8'hFF;
15'h3675:data=8'hFF;
15'h3676:data=8'hF8;
15'h3677:data=8'h00;
15'h3680:data=8'h00;
15'h3681:data=8'h00;
15'h3682:data=8'h03;
15'h3683:data=8'h0F;
15'h3684:data=8'h1F;
15'h3685:data=8'h3F;
15'h3686:data=8'h7E;
15'h3687:data=8'hF8;
15'h3688:data=8'hF0;
15'h3689:data=8'hF0;
15'h368a:data=8'hE0;
15'h368b:data=8'hE0;
15'h368c:data=8'hE0;
15'h368d:data=8'hE0;
15'h368e:data=8'hE0;
15'h368f:data=8'hF0;
15'h3690:data=8'hF0;
15'h3691:data=8'h7C;
15'h3692:data=8'h7F;
15'h3693:data=8'h3F;
15'h3694:data=8'h1F;
15'h3695:data=8'h07;
15'h3696:data=8'h00;
15'h3697:data=8'h00;
15'h36a0:data=8'h00;
15'h36a1:data=8'h00;
15'h36a2:data=8'h00;
15'h36a3:data=8'h00;
15'h36a4:data=8'h00;
15'h36a5:data=8'h00;
15'h36a6:data=8'h00;
15'h36a7:data=8'h00;
15'h36a8:data=8'h00;
15'h36a9:data=8'h00;
15'h36aa:data=8'h00;
15'h36ab:data=8'h00;
15'h36ac:data=8'h00;
15'h36ad:data=8'h00;
15'h36ae:data=8'h00;
15'h36af:data=8'h00;
15'h36b0:data=8'h00;
15'h36b1:data=8'h00;
15'h36b2:data=8'h00;
15'h36b3:data=8'h00;
15'h36b4:data=8'h00;
15'h36b5:data=8'h00;
15'h36b6:data=8'h00;
15'h36b7:data=8'h00;

15'h3700:data=8'h00;
15'h3701:data=8'h00;
15'h3702:data=8'h00;
15'h3703:data=8'h00;
15'h3704:data=8'h00;
15'h3705:data=8'h00;
15'h3706:data=8'h00;
15'h3707:data=8'h00;
15'h3708:data=8'h00;
15'h3709:data=8'h00;
15'h370a:data=8'h00;
15'h370b:data=8'h00;
15'h370c:data=8'h00;
15'h370d:data=8'h00;
15'h370e:data=8'h00;
15'h370f:data=8'h00;
15'h3710:data=8'h00;
15'h3711:data=8'h00;
15'h3712:data=8'h00;
15'h3713:data=8'h00;
15'h3714:data=8'h00;
15'h3715:data=8'h00;
15'h3716:data=8'h00;
15'h3717:data=8'h00;
15'h3720:data=8'h00;
15'h3721:data=8'h00;
15'h3722:data=8'h0F;
15'h3723:data=8'h0F;
15'h3724:data=8'h0F;
15'h3725:data=8'h0F;
15'h3726:data=8'h0F;
15'h3727:data=8'h0F;
15'h3728:data=8'h0F;
15'h3729:data=8'h0F;
15'h372a:data=8'h0F;
15'h372b:data=8'h0F;
15'h372c:data=8'h0F;
15'h372d:data=8'h0F;
15'h372e:data=8'h0F;
15'h372f:data=8'h0F;
15'h3730:data=8'hCF;
15'h3731:data=8'hEF;
15'h3732:data=8'hFF;
15'h3733:data=8'hFF;
15'h3734:data=8'h3F;
15'h3735:data=8'h0F;
15'h3736:data=8'h00;
15'h3737:data=8'h00;
15'h3740:data=8'h00;
15'h3741:data=8'h00;
15'h3742:data=8'h00;
15'h3743:data=8'h00;
15'h3744:data=8'h00;
15'h3745:data=8'h00;
15'h3746:data=8'h00;
15'h3747:data=8'h00;
15'h3748:data=8'h00;
15'h3749:data=8'h00;
15'h374a:data=8'h00;
15'h374b:data=8'h00;
15'h374c:data=8'hC0;
15'h374d:data=8'hF0;
15'h374e:data=8'hFC;
15'h374f:data=8'hFF;
15'h3750:data=8'h3F;
15'h3751:data=8'h0F;
15'h3752:data=8'h03;
15'h3753:data=8'h00;
15'h3754:data=8'h00;
15'h3755:data=8'h00;
15'h3756:data=8'h00;
15'h3757:data=8'h00;
15'h3760:data=8'h00;
15'h3761:data=8'h00;
15'h3762:data=8'h00;
15'h3763:data=8'h00;
15'h3764:data=8'h00;
15'h3765:data=8'h00;
15'h3766:data=8'h00;
15'h3767:data=8'h00;
15'h3768:data=8'h00;
15'h3769:data=8'hC0;
15'h376a:data=8'hF8;
15'h376b:data=8'hFE;
15'h376c:data=8'hFF;
15'h376d:data=8'h1F;
15'h376e:data=8'h03;
15'h376f:data=8'h00;
15'h3770:data=8'h00;
15'h3771:data=8'h00;
15'h3772:data=8'h00;
15'h3773:data=8'h00;
15'h3774:data=8'h00;
15'h3775:data=8'h00;
15'h3776:data=8'h00;
15'h3777:data=8'h00;
15'h3780:data=8'h00;
15'h3781:data=8'h00;
15'h3782:data=8'h00;
15'h3783:data=8'h00;
15'h3784:data=8'h00;
15'h3785:data=8'h00;
15'h3786:data=8'h80;
15'h3787:data=8'hF0;
15'h3788:data=8'hFF;
15'h3789:data=8'hFF;
15'h378a:data=8'hFF;
15'h378b:data=8'h0F;
15'h378c:data=8'h00;
15'h378d:data=8'h00;
15'h378e:data=8'h00;
15'h378f:data=8'h00;
15'h3790:data=8'h00;
15'h3791:data=8'h00;
15'h3792:data=8'h00;
15'h3793:data=8'h00;
15'h3794:data=8'h00;
15'h3795:data=8'h00;
15'h3796:data=8'h00;
15'h3797:data=8'h00;
15'h37a0:data=8'h00;
15'h37a1:data=8'h00;
15'h37a2:data=8'h00;
15'h37a3:data=8'h00;
15'h37a4:data=8'h00;
15'h37a5:data=8'h00;
15'h37a6:data=8'h00;
15'h37a7:data=8'h00;
15'h37a8:data=8'h00;
15'h37a9:data=8'h00;
15'h37aa:data=8'h00;
15'h37ab:data=8'h00;
15'h37ac:data=8'h00;
15'h37ad:data=8'h00;
15'h37ae:data=8'h00;
15'h37af:data=8'h00;
15'h37b0:data=8'h00;
15'h37b1:data=8'h00;
15'h37b2:data=8'h00;
15'h37b3:data=8'h00;
15'h37b4:data=8'h00;
15'h37b5:data=8'h00;
15'h37b6:data=8'h00;
15'h37b7:data=8'h00;

15'h3800:data=8'h00;
15'h3801:data=8'h00;
15'h3802:data=8'h00;
15'h3803:data=8'h00;
15'h3804:data=8'h00;
15'h3805:data=8'h00;
15'h3806:data=8'h00;
15'h3807:data=8'h00;
15'h3808:data=8'h00;
15'h3809:data=8'h00;
15'h380a:data=8'h00;
15'h380b:data=8'h00;
15'h380c:data=8'h00;
15'h380d:data=8'h00;
15'h380e:data=8'h00;
15'h380f:data=8'h00;
15'h3810:data=8'h00;
15'h3811:data=8'h00;
15'h3812:data=8'h00;
15'h3813:data=8'h00;
15'h3814:data=8'h00;
15'h3815:data=8'h00;
15'h3816:data=8'h00;
15'h3817:data=8'h00;
15'h3820:data=8'h00;
15'h3821:data=8'h00;
15'h3822:data=8'hC0;
15'h3823:data=8'hF0;
15'h3824:data=8'hFC;
15'h3825:data=8'hFE;
15'h3826:data=8'h1E;
15'h3827:data=8'h0F;
15'h3828:data=8'h07;
15'h3829:data=8'h07;
15'h382a:data=8'h07;
15'h382b:data=8'h07;
15'h382c:data=8'h07;
15'h382d:data=8'h07;
15'h382e:data=8'h0F;
15'h382f:data=8'h0F;
15'h3830:data=8'h3E;
15'h3831:data=8'hFE;
15'h3832:data=8'hFC;
15'h3833:data=8'hF8;
15'h3834:data=8'hC0;
15'h3835:data=8'h00;
15'h3836:data=8'h00;
15'h3837:data=8'h00;
15'h3840:data=8'h00;
15'h3841:data=8'h00;
15'h3842:data=8'h03;
15'h3843:data=8'h0F;
15'h3844:data=8'h3F;
15'h3845:data=8'hBF;
15'h3846:data=8'hFC;
15'h3847:data=8'hF0;
15'h3848:data=8'hE0;
15'h3849:data=8'hE0;
15'h384a:data=8'hE0;
15'h384b:data=8'hE0;
15'h384c:data=8'hE0;
15'h384d:data=8'hE0;
15'h384e:data=8'hF0;
15'h384f:data=8'hF8;
15'h3850:data=8'hFC;
15'h3851:data=8'h3F;
15'h3852:data=8'h1F;
15'h3853:data=8'h0F;
15'h3854:data=8'h01;
15'h3855:data=8'h00;
15'h3856:data=8'h00;
15'h3857:data=8'h00;
15'h3860:data=8'h00;
15'h3861:data=8'hE0;
15'h3862:data=8'hFC;
15'h3863:data=8'hFE;
15'h3864:data=8'hFF;
15'h3865:data=8'h1F;
15'h3866:data=8'h07;
15'h3867:data=8'h03;
15'h3868:data=8'h03;
15'h3869:data=8'h01;
15'h386a:data=8'h01;
15'h386b:data=8'h01;
15'h386c:data=8'h01;
15'h386d:data=8'h01;
15'h386e:data=8'h03;
15'h386f:data=8'h03;
15'h3870:data=8'h07;
15'h3871:data=8'h1F;
15'h3872:data=8'hFF;
15'h3873:data=8'hFE;
15'h3874:data=8'hFC;
15'h3875:data=8'hC0;
15'h3876:data=8'h00;
15'h3877:data=8'h00;
15'h3880:data=8'h00;
15'h3881:data=8'h01;
15'h3882:data=8'h0F;
15'h3883:data=8'h3F;
15'h3884:data=8'h7F;
15'h3885:data=8'h7E;
15'h3886:data=8'hF8;
15'h3887:data=8'hF0;
15'h3888:data=8'hF0;
15'h3889:data=8'hE0;
15'h388a:data=8'hE0;
15'h388b:data=8'hE0;
15'h388c:data=8'hE0;
15'h388d:data=8'hE0;
15'h388e:data=8'hF0;
15'h388f:data=8'hF0;
15'h3890:data=8'hF8;
15'h3891:data=8'h7E;
15'h3892:data=8'h3F;
15'h3893:data=8'h1F;
15'h3894:data=8'h0F;
15'h3895:data=8'h00;
15'h3896:data=8'h00;
15'h3897:data=8'h00;
15'h38a0:data=8'h00;
15'h38a1:data=8'h00;
15'h38a2:data=8'h00;
15'h38a3:data=8'h00;
15'h38a4:data=8'h00;
15'h38a5:data=8'h00;
15'h38a6:data=8'h00;
15'h38a7:data=8'h00;
15'h38a8:data=8'h00;
15'h38a9:data=8'h00;
15'h38aa:data=8'h00;
15'h38ab:data=8'h00;
15'h38ac:data=8'h00;
15'h38ad:data=8'h00;
15'h38ae:data=8'h00;
15'h38af:data=8'h00;
15'h38b0:data=8'h00;
15'h38b1:data=8'h00;
15'h38b2:data=8'h00;
15'h38b3:data=8'h00;
15'h38b4:data=8'h00;
15'h38b5:data=8'h00;
15'h38b6:data=8'h00;
15'h38b7:data=8'h00;

15'h3900:data=8'h00;
15'h3901:data=8'h00;
15'h3902:data=8'h00;
15'h3903:data=8'h00;
15'h3904:data=8'h00;
15'h3905:data=8'h00;
15'h3906:data=8'h00;
15'h3907:data=8'h00;
15'h3908:data=8'h00;
15'h3909:data=8'h00;
15'h390a:data=8'h80;
15'h390b:data=8'h80;
15'h390c:data=8'h80;
15'h390d:data=8'h00;
15'h390e:data=8'h00;
15'h390f:data=8'h00;
15'h3910:data=8'h00;
15'h3911:data=8'h00;
15'h3912:data=8'h00;
15'h3913:data=8'h00;
15'h3914:data=8'h00;
15'h3915:data=8'h00;
15'h3916:data=8'h00;
15'h3917:data=8'h00;
15'h3920:data=8'h00;
15'h3921:data=8'h80;
15'h3922:data=8'hF0;
15'h3923:data=8'hF8;
15'h3924:data=8'hFC;
15'h3925:data=8'h7E;
15'h3926:data=8'h1E;
15'h3927:data=8'h0F;
15'h3928:data=8'h0F;
15'h3929:data=8'h07;
15'h392a:data=8'h07;
15'h392b:data=8'h07;
15'h392c:data=8'h07;
15'h392d:data=8'h0F;
15'h392e:data=8'h0F;
15'h392f:data=8'h1F;
15'h3930:data=8'h7E;
15'h3931:data=8'hFC;
15'h3932:data=8'hFC;
15'h3933:data=8'hF0;
15'h3934:data=8'hE0;
15'h3935:data=8'h00;
15'h3936:data=8'h00;
15'h3937:data=8'h00;
15'h3940:data=8'h00;
15'h3941:data=8'h3F;
15'h3942:data=8'hFF;
15'h3943:data=8'hFF;
15'h3944:data=8'hFF;
15'h3945:data=8'hE0;
15'h3946:data=8'h80;
15'h3947:data=8'h00;
15'h3948:data=8'h00;
15'h3949:data=8'h00;
15'h394a:data=8'h00;
15'h394b:data=8'h00;
15'h394c:data=8'h00;
15'h394d:data=8'h00;
15'h394e:data=8'h80;
15'h394f:data=8'hC0;
15'h3950:data=8'hE0;
15'h3951:data=8'hFF;
15'h3952:data=8'hFF;
15'h3953:data=8'hFF;
15'h3954:data=8'h1F;
15'h3955:data=8'h00;
15'h3956:data=8'h00;
15'h3957:data=8'h00;
15'h3960:data=8'h00;
15'h3961:data=8'h00;
15'h3962:data=8'h00;
15'h3963:data=8'h03;
15'h3964:data=8'h03;
15'h3965:data=8'h07;
15'h3966:data=8'h07;
15'h3967:data=8'h0F;
15'h3968:data=8'h0F;
15'h3969:data=8'h0E;
15'h396a:data=8'h0E;
15'h396b:data=8'hCE;
15'h396c:data=8'hFE;
15'h396d:data=8'hFF;
15'h396e:data=8'hFF;
15'h396f:data=8'h7F;
15'h3970:data=8'h1F;
15'h3971:data=8'h0F;
15'h3972:data=8'h03;
15'h3973:data=8'h00;
15'h3974:data=8'h00;
15'h3975:data=8'h00;
15'h3976:data=8'h00;
15'h3977:data=8'h00;
15'h3980:data=8'h00;
15'h3981:data=8'h00;
15'h3982:data=8'h00;
15'h3983:data=8'h00;
15'h3984:data=8'h00;
15'h3985:data=8'h00;
15'h3986:data=8'h00;
15'h3987:data=8'hC0;
15'h3988:data=8'hF0;
15'h3989:data=8'hFC;
15'h398a:data=8'hFF;
15'h398b:data=8'h3F;
15'h398c:data=8'h0F;
15'h398d:data=8'h07;
15'h398e:data=8'h01;
15'h398f:data=8'h00;
15'h3990:data=8'h00;
15'h3991:data=8'h00;
15'h3992:data=8'h00;
15'h3993:data=8'h00;
15'h3994:data=8'h00;
15'h3995:data=8'h00;
15'h3996:data=8'h00;
15'h3997:data=8'h00;
15'h39a0:data=8'h00;
15'h39a1:data=8'h00;
15'h39a2:data=8'h00;
15'h39a3:data=8'h00;
15'h39a4:data=8'h00;
15'h39a5:data=8'h00;
15'h39a6:data=8'h00;
15'h39a7:data=8'h00;
15'h39a8:data=8'h00;
15'h39a9:data=8'h00;
15'h39aa:data=8'h00;
15'h39ab:data=8'h00;
15'h39ac:data=8'h00;
15'h39ad:data=8'h00;
15'h39ae:data=8'h00;
15'h39af:data=8'h00;
15'h39b0:data=8'h00;
15'h39b1:data=8'h00;
15'h39b2:data=8'h00;
15'h39b3:data=8'h00;
15'h39b4:data=8'h00;
15'h39b5:data=8'h00;
15'h39b6:data=8'h00;
15'h39b7:data=8'h00;


		default:data=8'h00;
		endcase
	end
	
endmodule
