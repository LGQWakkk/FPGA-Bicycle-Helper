`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/06/15 16:17:11
// Design Name: 
// Module Name: pic_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pic_rom(
	input wire clk,
	input wire [13:0] addr,
	output reg [7:0] data
    );
	
	reg [13:0] addr_reg;
	
	always@(posedge clk)begin
		addr_reg<=addr;
	end
	
	always@(*)begin
		case(addr_reg)
		/////////////////////////////////////////////////////////PIC1 Speed
14'h0000:data=8'h00;
14'h0001:data=8'h00;
14'h0002:data=8'h00;
14'h0003:data=8'h00;
14'h0004:data=8'h00;
14'h0005:data=8'h00;
14'h0006:data=8'h00;
14'h0007:data=8'h00;
14'h0008:data=8'h00;
14'h0009:data=8'h00;
14'h000a:data=8'h00;
14'h000b:data=8'h00;
14'h000c:data=8'h00;
14'h000d:data=8'h00;
14'h000e:data=8'h00;
14'h000f:data=8'h00;
14'h0010:data=8'h00;
14'h0011:data=8'h00;
14'h0012:data=8'h00;
14'h0013:data=8'h00;
14'h0014:data=8'h00;
14'h0015:data=8'h00;
14'h0016:data=8'h00;
14'h0017:data=8'h00;
14'h0018:data=8'h00;
14'h0019:data=8'h00;
14'h001a:data=8'h00;
14'h001b:data=8'h00;
14'h001c:data=8'h00;
14'h001d:data=8'h00;
14'h001e:data=8'h00;
14'h001f:data=8'h00;
14'h0020:data=8'h00;
14'h0021:data=8'h00;
14'h0022:data=8'h00;
14'h0023:data=8'h00;
14'h0024:data=8'h00;
14'h0025:data=8'h00;
14'h0026:data=8'h00;
14'h0027:data=8'h00;
14'h0028:data=8'h00;
14'h0029:data=8'h00;
14'h002a:data=8'h00;
14'h002b:data=8'h00;
14'h002c:data=8'h00;
14'h002d:data=8'h00;
14'h002e:data=8'h00;
14'h002f:data=8'h00;
14'h0030:data=8'h00;
14'h0031:data=8'h00;
14'h0032:data=8'h00;
14'h0033:data=8'h00;
14'h0034:data=8'h00;
14'h0035:data=8'h00;
14'h0036:data=8'h00;
14'h0037:data=8'h00;
14'h0038:data=8'h00;
14'h0039:data=8'h00;
14'h003a:data=8'h00;
14'h003b:data=8'h00;
14'h003c:data=8'h00;
14'h003d:data=8'h00;
14'h003e:data=8'h00;
14'h003f:data=8'h00;
14'h0040:data=8'h00;
14'h0041:data=8'h00;
14'h0042:data=8'h00;
14'h0043:data=8'h00;
14'h0044:data=8'h00;
14'h0045:data=8'h00;
14'h0046:data=8'h00;
14'h0047:data=8'h00;
14'h0048:data=8'h00;
14'h0049:data=8'h00;
14'h004a:data=8'h00;
14'h004b:data=8'h00;
14'h004c:data=8'h00;
14'h004d:data=8'h00;
14'h004e:data=8'h00;
14'h004f:data=8'h00;
14'h0050:data=8'h00;
14'h0051:data=8'h00;
14'h0052:data=8'h00;
14'h0053:data=8'h00;
14'h0054:data=8'h00;
14'h0055:data=8'h00;
14'h0056:data=8'h00;
14'h0057:data=8'h00;
14'h0058:data=8'h00;
14'h0059:data=8'h00;
14'h005a:data=8'h00;
14'h005b:data=8'h00;
14'h005c:data=8'h00;
14'h005d:data=8'h00;
14'h005e:data=8'h00;
14'h005f:data=8'h00;
14'h0060:data=8'h00;
14'h0061:data=8'h00;
14'h0062:data=8'h00;
14'h0063:data=8'h00;
14'h0064:data=8'h00;
14'h0065:data=8'h00;
14'h0066:data=8'h00;
14'h0067:data=8'h00;
14'h0068:data=8'h00;
14'h0069:data=8'h00;
14'h006a:data=8'h00;
14'h006b:data=8'h00;
14'h006c:data=8'h00;
14'h006d:data=8'h00;
14'h006e:data=8'h00;
14'h006f:data=8'h00;
14'h0070:data=8'h00;
14'h0071:data=8'h00;
14'h0072:data=8'h00;
14'h0073:data=8'h00;
14'h0074:data=8'h00;
14'h0075:data=8'h00;
14'h0076:data=8'h00;
14'h0077:data=8'h00;
14'h0078:data=8'h00;
14'h0079:data=8'h00;
14'h007a:data=8'h00;
14'h007b:data=8'h00;
14'h007c:data=8'h00;
14'h007d:data=8'h00;
14'h007e:data=8'h00;
14'h007f:data=8'h00;
14'h0800:data=8'h00;
14'h0801:data=8'h00;
14'h0802:data=8'h00;
14'h0803:data=8'h00;
14'h0804:data=8'h00;
14'h0805:data=8'h00;
14'h0806:data=8'h00;
14'h0807:data=8'h00;
14'h0808:data=8'h00;
14'h0809:data=8'h00;
14'h080a:data=8'h80;
14'h080b:data=8'h80;
14'h080c:data=8'hC0;
14'h080d:data=8'hC0;
14'h080e:data=8'hE0;
14'h080f:data=8'hE0;
14'h0810:data=8'hE0;
14'h0811:data=8'hE0;
14'h0812:data=8'hE0;
14'h0813:data=8'hE0;
14'h0814:data=8'hE0;
14'h0815:data=8'hE0;
14'h0816:data=8'hE0;
14'h0817:data=8'hE0;
14'h0818:data=8'hE0;
14'h0819:data=8'hC0;
14'h081a:data=8'hC0;
14'h081b:data=8'h80;
14'h081c:data=8'h00;
14'h081d:data=8'h00;
14'h081e:data=8'h00;
14'h081f:data=8'h00;
14'h0820:data=8'h00;
14'h0821:data=8'h00;
14'h0822:data=8'h00;
14'h0823:data=8'h00;
14'h0824:data=8'h00;
14'h0825:data=8'h00;
14'h0826:data=8'h00;
14'h0827:data=8'h00;
14'h0828:data=8'h00;
14'h0829:data=8'h00;
14'h082a:data=8'h00;
14'h082b:data=8'h00;
14'h082c:data=8'h00;
14'h082d:data=8'h00;
14'h082e:data=8'h00;
14'h082f:data=8'h00;
14'h0830:data=8'h00;
14'h0831:data=8'h00;
14'h0832:data=8'h00;
14'h0833:data=8'h00;
14'h0834:data=8'h00;
14'h0835:data=8'h00;
14'h0836:data=8'h00;
14'h0837:data=8'h00;
14'h0838:data=8'h00;
14'h0839:data=8'h00;
14'h083a:data=8'h00;
14'h083b:data=8'h00;
14'h083c:data=8'h00;
14'h083d:data=8'h00;
14'h083e:data=8'h00;
14'h083f:data=8'h00;
14'h0840:data=8'h00;
14'h0841:data=8'h00;
14'h0842:data=8'h00;
14'h0843:data=8'h00;
14'h0844:data=8'h00;
14'h0845:data=8'h00;
14'h0846:data=8'h00;
14'h0847:data=8'h00;
14'h0848:data=8'h00;
14'h0849:data=8'h00;
14'h084a:data=8'h00;
14'h084b:data=8'h00;
14'h084c:data=8'h00;
14'h084d:data=8'h00;
14'h084e:data=8'h00;
14'h084f:data=8'h00;
14'h0850:data=8'h00;
14'h0851:data=8'h00;
14'h0852:data=8'h00;
14'h0853:data=8'h00;
14'h0854:data=8'h00;
14'h0855:data=8'h00;
14'h0856:data=8'h00;
14'h0857:data=8'h00;
14'h0858:data=8'h00;
14'h0859:data=8'h00;
14'h085a:data=8'h00;
14'h085b:data=8'h00;
14'h085c:data=8'h00;
14'h085d:data=8'h00;
14'h085e:data=8'h00;
14'h085f:data=8'h00;
14'h0860:data=8'h00;
14'h0861:data=8'h00;
14'h0862:data=8'h00;
14'h0863:data=8'h00;
14'h0864:data=8'h00;
14'h0865:data=8'h00;
14'h0866:data=8'h00;
14'h0867:data=8'h00;
14'h0868:data=8'h00;
14'h0869:data=8'h00;
14'h086a:data=8'h00;
14'h086b:data=8'h00;
14'h086c:data=8'h00;
14'h086d:data=8'h00;
14'h086e:data=8'h00;
14'h086f:data=8'h00;
14'h0870:data=8'h00;
14'h0871:data=8'h00;
14'h0872:data=8'hE0;
14'h0873:data=8'hF0;
14'h0874:data=8'hF0;
14'h0875:data=8'hF0;
14'h0876:data=8'hF0;
14'h0877:data=8'hF0;
14'h0878:data=8'hF0;
14'h0879:data=8'hF0;
14'h087a:data=8'hF0;
14'h087b:data=8'h00;
14'h087c:data=8'h00;
14'h087d:data=8'h00;
14'h087e:data=8'h00;
14'h087f:data=8'h00;
14'h1000:data=8'h00;
14'h1001:data=8'h00;
14'h1002:data=8'h00;
14'h1003:data=8'h00;
14'h1004:data=8'h00;
14'h1005:data=8'h00;
14'h1006:data=8'h00;
14'h1007:data=8'hE0;
14'h1008:data=8'hFC;
14'h1009:data=8'hFF;
14'h100a:data=8'hFF;
14'h100b:data=8'hFF;
14'h100c:data=8'hFF;
14'h100d:data=8'hFF;
14'h100e:data=8'hFF;
14'h100f:data=8'hFF;
14'h1010:data=8'hBF;
14'h1011:data=8'h1F;
14'h1012:data=8'h1F;
14'h1013:data=8'h0F;
14'h1014:data=8'h1F;
14'h1015:data=8'h1F;
14'h1016:data=8'h1F;
14'h1017:data=8'h1F;
14'h1018:data=8'h3F;
14'h1019:data=8'h3F;
14'h101a:data=8'h3F;
14'h101b:data=8'h1F;
14'h101c:data=8'h00;
14'h101d:data=8'h00;
14'h101e:data=8'hE0;
14'h101f:data=8'hE0;
14'h1020:data=8'hE0;
14'h1021:data=8'hE0;
14'h1022:data=8'hE0;
14'h1023:data=8'hE0;
14'h1024:data=8'hE0;
14'h1025:data=8'hE0;
14'h1026:data=8'hC0;
14'h1027:data=8'hE0;
14'h1028:data=8'hE0;
14'h1029:data=8'hE0;
14'h102a:data=8'hE0;
14'h102b:data=8'hE0;
14'h102c:data=8'hE0;
14'h102d:data=8'hE0;
14'h102e:data=8'hE0;
14'h102f:data=8'hC0;
14'h1030:data=8'hC0;
14'h1031:data=8'h80;
14'h1032:data=8'h00;
14'h1033:data=8'h00;
14'h1034:data=8'h00;
14'h1035:data=8'h00;
14'h1036:data=8'h00;
14'h1037:data=8'h00;
14'h1038:data=8'h00;
14'h1039:data=8'h80;
14'h103a:data=8'h80;
14'h103b:data=8'hC0;
14'h103c:data=8'hC0;
14'h103d:data=8'hE0;
14'h103e:data=8'hE0;
14'h103f:data=8'hE0;
14'h1040:data=8'hE0;
14'h1041:data=8'hE0;
14'h1042:data=8'hE0;
14'h1043:data=8'hE0;
14'h1044:data=8'hE0;
14'h1045:data=8'hE0;
14'h1046:data=8'hC0;
14'h1047:data=8'hC0;
14'h1048:data=8'h80;
14'h1049:data=8'h00;
14'h104a:data=8'h00;
14'h104b:data=8'h00;
14'h104c:data=8'h00;
14'h104d:data=8'h00;
14'h104e:data=8'h00;
14'h104f:data=8'h80;
14'h1050:data=8'hC0;
14'h1051:data=8'hC0;
14'h1052:data=8'hE0;
14'h1053:data=8'hE0;
14'h1054:data=8'hE0;
14'h1055:data=8'hE0;
14'h1056:data=8'hE0;
14'h1057:data=8'hE0;
14'h1058:data=8'hE0;
14'h1059:data=8'hE0;
14'h105a:data=8'hE0;
14'h105b:data=8'hE0;
14'h105c:data=8'hC0;
14'h105d:data=8'hC0;
14'h105e:data=8'h80;
14'h105f:data=8'h00;
14'h1060:data=8'h00;
14'h1061:data=8'h00;
14'h1062:data=8'h00;
14'h1063:data=8'h00;
14'h1064:data=8'h00;
14'h1065:data=8'h80;
14'h1066:data=8'h80;
14'h1067:data=8'hC0;
14'h1068:data=8'hC0;
14'h1069:data=8'hE0;
14'h106a:data=8'hE0;
14'h106b:data=8'hE0;
14'h106c:data=8'hE0;
14'h106d:data=8'hE0;
14'h106e:data=8'hE0;
14'h106f:data=8'hE0;
14'h1070:data=8'hE0;
14'h1071:data=8'hFC;
14'h1072:data=8'hFF;
14'h1073:data=8'hFF;
14'h1074:data=8'hFF;
14'h1075:data=8'hFF;
14'h1076:data=8'hFF;
14'h1077:data=8'hFF;
14'h1078:data=8'hFF;
14'h1079:data=8'h1F;
14'h107a:data=8'h00;
14'h107b:data=8'h00;
14'h107c:data=8'h00;
14'h107d:data=8'h00;
14'h107e:data=8'h00;
14'h107f:data=8'h00;
14'h1800:data=8'h00;
14'h1801:data=8'h00;
14'h1802:data=8'h00;
14'h1803:data=8'h00;
14'h1804:data=8'h00;
14'h1805:data=8'h00;
14'h1806:data=8'h00;
14'h1807:data=8'h01;
14'h1808:data=8'h0F;
14'h1809:data=8'h3F;
14'h180a:data=8'h7F;
14'h180b:data=8'hFF;
14'h180c:data=8'hFF;
14'h180d:data=8'hFF;
14'h180e:data=8'hFF;
14'h180f:data=8'hFF;
14'h1810:data=8'hFF;
14'h1811:data=8'hFF;
14'h1812:data=8'hFE;
14'h1813:data=8'hFC;
14'h1814:data=8'hFC;
14'h1815:data=8'hF8;
14'h1816:data=8'hF0;
14'h1817:data=8'hE0;
14'h1818:data=8'hC0;
14'h1819:data=8'h00;
14'h181a:data=8'h00;
14'h181b:data=8'h00;
14'h181c:data=8'h00;
14'h181d:data=8'hF8;
14'h181e:data=8'hFF;
14'h181f:data=8'hFF;
14'h1820:data=8'hFF;
14'h1821:data=8'hFF;
14'h1822:data=8'hFF;
14'h1823:data=8'hFF;
14'h1824:data=8'hFF;
14'h1825:data=8'hFF;
14'h1826:data=8'h7F;
14'h1827:data=8'h3F;
14'h1828:data=8'h1F;
14'h1829:data=8'h1F;
14'h182a:data=8'h1F;
14'h182b:data=8'hFF;
14'h182c:data=8'hFF;
14'h182d:data=8'hFF;
14'h182e:data=8'hFF;
14'h182f:data=8'hFF;
14'h1830:data=8'hFF;
14'h1831:data=8'hFF;
14'h1832:data=8'hFE;
14'h1833:data=8'hE0;
14'h1834:data=8'h00;
14'h1835:data=8'hF0;
14'h1836:data=8'hFC;
14'h1837:data=8'hFE;
14'h1838:data=8'hFF;
14'h1839:data=8'hFF;
14'h183a:data=8'hFF;
14'h183b:data=8'hFF;
14'h183c:data=8'hFF;
14'h183d:data=8'hFF;
14'h183e:data=8'hFF;
14'h183f:data=8'hEF;
14'h1840:data=8'hEF;
14'h1841:data=8'hFF;
14'h1842:data=8'hFF;
14'h1843:data=8'hFF;
14'h1844:data=8'hFF;
14'h1845:data=8'hFF;
14'h1846:data=8'hFF;
14'h1847:data=8'hFF;
14'h1848:data=8'hFF;
14'h1849:data=8'hFF;
14'h184a:data=8'h80;
14'h184b:data=8'hF0;
14'h184c:data=8'hFC;
14'h184d:data=8'hFE;
14'h184e:data=8'hFF;
14'h184f:data=8'hFF;
14'h1850:data=8'hFF;
14'h1851:data=8'hFF;
14'h1852:data=8'hFF;
14'h1853:data=8'hFF;
14'h1854:data=8'hFF;
14'h1855:data=8'hEF;
14'h1856:data=8'hEF;
14'h1857:data=8'hFF;
14'h1858:data=8'hFF;
14'h1859:data=8'hFF;
14'h185a:data=8'hFF;
14'h185b:data=8'hFF;
14'h185c:data=8'hFF;
14'h185d:data=8'hFF;
14'h185e:data=8'hFF;
14'h185f:data=8'hFE;
14'h1860:data=8'h80;
14'h1861:data=8'hF0;
14'h1862:data=8'hFC;
14'h1863:data=8'hFE;
14'h1864:data=8'hFF;
14'h1865:data=8'hFF;
14'h1866:data=8'hFF;
14'h1867:data=8'hFF;
14'h1868:data=8'hFF;
14'h1869:data=8'hFF;
14'h186a:data=8'h7F;
14'h186b:data=8'h3F;
14'h186c:data=8'h1F;
14'h186d:data=8'h1F;
14'h186e:data=8'h0F;
14'h186f:data=8'hFF;
14'h1870:data=8'hFF;
14'h1871:data=8'hFF;
14'h1872:data=8'hFF;
14'h1873:data=8'hFF;
14'h1874:data=8'hFF;
14'h1875:data=8'hFF;
14'h1876:data=8'hFF;
14'h1877:data=8'h7F;
14'h1878:data=8'h03;
14'h1879:data=8'h00;
14'h187a:data=8'h00;
14'h187b:data=8'h00;
14'h187c:data=8'h00;
14'h187d:data=8'h00;
14'h187e:data=8'h00;
14'h187f:data=8'h00;
14'h2000:data=8'h00;
14'h2001:data=8'h00;
14'h2002:data=8'h00;
14'h2003:data=8'h00;
14'h2004:data=8'h80;
14'h2005:data=8'hF8;
14'h2006:data=8'hF8;
14'h2007:data=8'hF0;
14'h2008:data=8'hF0;
14'h2009:data=8'hE0;
14'h200a:data=8'hE0;
14'h200b:data=8'hE0;
14'h200c:data=8'hC0;
14'h200d:data=8'hC1;
14'h200e:data=8'hE1;
14'h200f:data=8'hE3;
14'h2010:data=8'hF7;
14'h2011:data=8'hFF;
14'h2012:data=8'hFF;
14'h2013:data=8'hFF;
14'h2014:data=8'hFF;
14'h2015:data=8'hFF;
14'h2016:data=8'hFF;
14'h2017:data=8'hFF;
14'h2018:data=8'hFF;
14'h2019:data=8'h7F;
14'h201a:data=8'h00;
14'h201b:data=8'hE0;
14'h201c:data=8'hFF;
14'h201d:data=8'hFF;
14'h201e:data=8'hFF;
14'h201f:data=8'hFF;
14'h2020:data=8'hFF;
14'h2021:data=8'hFF;
14'h2022:data=8'hFF;
14'h2023:data=8'hFF;
14'h2024:data=8'hCF;
14'h2025:data=8'hC1;
14'h2026:data=8'hE0;
14'h2027:data=8'hE0;
14'h2028:data=8'hF0;
14'h2029:data=8'hF8;
14'h202a:data=8'hFE;
14'h202b:data=8'hFF;
14'h202c:data=8'hFF;
14'h202d:data=8'hFF;
14'h202e:data=8'hFF;
14'h202f:data=8'hFF;
14'h2030:data=8'hFF;
14'h2031:data=8'h7F;
14'h2032:data=8'h1F;
14'h2033:data=8'h00;
14'h2034:data=8'h3F;
14'h2035:data=8'hFF;
14'h2036:data=8'hFF;
14'h2037:data=8'hFF;
14'h2038:data=8'hFF;
14'h2039:data=8'hFF;
14'h203a:data=8'hFF;
14'h203b:data=8'hFF;
14'h203c:data=8'hFF;
14'h203d:data=8'hEF;
14'h203e:data=8'hCF;
14'h203f:data=8'hCF;
14'h2040:data=8'hEF;
14'h2041:data=8'hEF;
14'h2042:data=8'hEF;
14'h2043:data=8'hEF;
14'h2044:data=8'hF7;
14'h2045:data=8'hF7;
14'h2046:data=8'hFF;
14'h2047:data=8'h73;
14'h2048:data=8'h03;
14'h2049:data=8'h00;
14'h204a:data=8'hFF;
14'h204b:data=8'hFF;
14'h204c:data=8'hFF;
14'h204d:data=8'hFF;
14'h204e:data=8'hFF;
14'h204f:data=8'hFF;
14'h2050:data=8'hFF;
14'h2051:data=8'hFF;
14'h2052:data=8'hFF;
14'h2053:data=8'hEF;
14'h2054:data=8'hCF;
14'h2055:data=8'hCF;
14'h2056:data=8'hEF;
14'h2057:data=8'hEF;
14'h2058:data=8'hEF;
14'h2059:data=8'hEF;
14'h205a:data=8'hF7;
14'h205b:data=8'hFF;
14'h205c:data=8'hF7;
14'h205d:data=8'h03;
14'h205e:data=8'h01;
14'h205f:data=8'h00;
14'h2060:data=8'hFF;
14'h2061:data=8'hFF;
14'h2062:data=8'hFF;
14'h2063:data=8'hFF;
14'h2064:data=8'hFF;
14'h2065:data=8'hFF;
14'h2066:data=8'hFF;
14'h2067:data=8'hFF;
14'h2068:data=8'hFF;
14'h2069:data=8'hC0;
14'h206a:data=8'hE0;
14'h206b:data=8'hE0;
14'h206c:data=8'hF0;
14'h206d:data=8'hFC;
14'h206e:data=8'hFF;
14'h206f:data=8'hFF;
14'h2070:data=8'hFF;
14'h2071:data=8'hFF;
14'h2072:data=8'hFF;
14'h2073:data=8'hFF;
14'h2074:data=8'hFF;
14'h2075:data=8'hFF;
14'h2076:data=8'h0F;
14'h2077:data=8'h00;
14'h2078:data=8'h00;
14'h2079:data=8'h00;
14'h207a:data=8'h00;
14'h207b:data=8'h00;
14'h207c:data=8'h00;
14'h207d:data=8'h00;
14'h207e:data=8'h00;
14'h207f:data=8'h00;
14'h2800:data=8'h00;
14'h2801:data=8'h00;
14'h2802:data=8'h00;
14'h2803:data=8'h00;
14'h2804:data=8'h07;
14'h2805:data=8'h0F;
14'h2806:data=8'h0F;
14'h2807:data=8'h1F;
14'h2808:data=8'h1F;
14'h2809:data=8'h1F;
14'h280a:data=8'h1F;
14'h280b:data=8'h1F;
14'h280c:data=8'h1F;
14'h280d:data=8'h1F;
14'h280e:data=8'h1F;
14'h280f:data=8'h1F;
14'h2810:data=8'h1F;
14'h2811:data=8'h1F;
14'h2812:data=8'h1F;
14'h2813:data=8'h1F;
14'h2814:data=8'h0F;
14'h2815:data=8'h0F;
14'h2816:data=8'h07;
14'h2817:data=8'h07;
14'h2818:data=8'h01;
14'h2819:data=8'h80;
14'h281a:data=8'hFC;
14'h281b:data=8'hFF;
14'h281c:data=8'hFF;
14'h281d:data=8'hFF;
14'h281e:data=8'hFF;
14'h281f:data=8'hFF;
14'h2820:data=8'hFF;
14'h2821:data=8'hFF;
14'h2822:data=8'h3F;
14'h2823:data=8'h1F;
14'h2824:data=8'h1F;
14'h2825:data=8'h1F;
14'h2826:data=8'h1F;
14'h2827:data=8'h1F;
14'h2828:data=8'h1F;
14'h2829:data=8'h1F;
14'h282a:data=8'h1F;
14'h282b:data=8'h0F;
14'h282c:data=8'h0F;
14'h282d:data=8'h07;
14'h282e:data=8'h07;
14'h282f:data=8'h03;
14'h2830:data=8'h01;
14'h2831:data=8'h00;
14'h2832:data=8'h00;
14'h2833:data=8'h00;
14'h2834:data=8'h00;
14'h2835:data=8'h01;
14'h2836:data=8'h07;
14'h2837:data=8'h0F;
14'h2838:data=8'h0F;
14'h2839:data=8'h1F;
14'h283a:data=8'h1F;
14'h283b:data=8'h1F;
14'h283c:data=8'h1F;
14'h283d:data=8'h1F;
14'h283e:data=8'h1F;
14'h283f:data=8'h1F;
14'h2840:data=8'h1F;
14'h2841:data=8'h1F;
14'h2842:data=8'h1F;
14'h2843:data=8'h1F;
14'h2844:data=8'h0F;
14'h2845:data=8'h0F;
14'h2846:data=8'h0F;
14'h2847:data=8'h00;
14'h2848:data=8'h00;
14'h2849:data=8'h00;
14'h284a:data=8'h00;
14'h284b:data=8'h03;
14'h284c:data=8'h07;
14'h284d:data=8'h0F;
14'h284e:data=8'h0F;
14'h284f:data=8'h1F;
14'h2850:data=8'h1F;
14'h2851:data=8'h1F;
14'h2852:data=8'h1F;
14'h2853:data=8'h1F;
14'h2854:data=8'h1F;
14'h2855:data=8'h1F;
14'h2856:data=8'h1F;
14'h2857:data=8'h1F;
14'h2858:data=8'h1F;
14'h2859:data=8'h1F;
14'h285a:data=8'h0F;
14'h285b:data=8'h0F;
14'h285c:data=8'h07;
14'h285d:data=8'h00;
14'h285e:data=8'h00;
14'h285f:data=8'h00;
14'h2860:data=8'h01;
14'h2861:data=8'h07;
14'h2862:data=8'h0F;
14'h2863:data=8'h1F;
14'h2864:data=8'h1F;
14'h2865:data=8'h1F;
14'h2866:data=8'h1F;
14'h2867:data=8'h1F;
14'h2868:data=8'h1F;
14'h2869:data=8'h1F;
14'h286a:data=8'h1F;
14'h286b:data=8'h1F;
14'h286c:data=8'h0F;
14'h286d:data=8'h1F;
14'h286e:data=8'h1F;
14'h286f:data=8'h1F;
14'h2870:data=8'h1F;
14'h2871:data=8'h1F;
14'h2872:data=8'h1F;
14'h2873:data=8'h1F;
14'h2874:data=8'h1F;
14'h2875:data=8'h03;
14'h2876:data=8'h00;
14'h2877:data=8'h00;
14'h2878:data=8'h00;
14'h2879:data=8'h00;
14'h287a:data=8'h00;
14'h287b:data=8'h00;
14'h287c:data=8'h00;
14'h287d:data=8'h00;
14'h287e:data=8'h00;
14'h287f:data=8'h00;
14'h3000:data=8'h00;
14'h3001:data=8'h00;
14'h3002:data=8'h00;
14'h3003:data=8'h00;
14'h3004:data=8'h00;
14'h3005:data=8'h00;
14'h3006:data=8'h00;
14'h3007:data=8'h00;
14'h3008:data=8'h00;
14'h3009:data=8'h00;
14'h300a:data=8'h00;
14'h300b:data=8'h00;
14'h300c:data=8'h00;
14'h300d:data=8'h00;
14'h300e:data=8'h00;
14'h300f:data=8'h00;
14'h3010:data=8'h00;
14'h3011:data=8'h00;
14'h3012:data=8'h00;
14'h3013:data=8'h00;
14'h3014:data=8'h00;
14'h3015:data=8'h00;
14'h3016:data=8'h00;
14'h3017:data=8'h00;
14'h3018:data=8'h70;
14'h3019:data=8'h7F;
14'h301a:data=8'h7F;
14'h301b:data=8'h7F;
14'h301c:data=8'h7F;
14'h301d:data=8'h7F;
14'h301e:data=8'h7F;
14'h301f:data=8'h7F;
14'h3020:data=8'h7F;
14'h3021:data=8'h07;
14'h3022:data=8'h00;
14'h3023:data=8'h00;
14'h3024:data=8'h00;
14'h3025:data=8'h00;
14'h3026:data=8'h00;
14'h3027:data=8'h00;
14'h3028:data=8'h00;
14'h3029:data=8'h00;
14'h302a:data=8'h00;
14'h302b:data=8'h04;
14'h302c:data=8'h04;
14'h302d:data=8'h04;
14'h302e:data=8'h04;
14'h302f:data=8'h14;
14'h3030:data=8'h14;
14'h3031:data=8'h14;
14'h3032:data=8'h14;
14'h3033:data=8'h54;
14'h3034:data=8'h54;
14'h3035:data=8'h54;
14'h3036:data=8'h54;
14'h3037:data=8'h54;
14'h3038:data=8'h54;
14'h3039:data=8'h54;
14'h303a:data=8'h54;
14'h303b:data=8'h54;
14'h303c:data=8'h54;
14'h303d:data=8'h54;
14'h303e:data=8'h54;
14'h303f:data=8'h54;
14'h3040:data=8'h54;
14'h3041:data=8'h54;
14'h3042:data=8'h54;
14'h3043:data=8'h54;
14'h3044:data=8'h54;
14'h3045:data=8'h54;
14'h3046:data=8'h54;
14'h3047:data=8'h54;
14'h3048:data=8'h54;
14'h3049:data=8'h54;
14'h304a:data=8'h54;
14'h304b:data=8'h54;
14'h304c:data=8'h54;
14'h304d:data=8'h54;
14'h304e:data=8'h54;
14'h304f:data=8'h54;
14'h3050:data=8'h54;
14'h3051:data=8'h54;
14'h3052:data=8'h54;
14'h3053:data=8'h54;
14'h3054:data=8'h54;
14'h3055:data=8'h54;
14'h3056:data=8'h54;
14'h3057:data=8'h54;
14'h3058:data=8'h54;
14'h3059:data=8'h54;
14'h305a:data=8'h54;
14'h305b:data=8'h54;
14'h305c:data=8'h54;
14'h305d:data=8'h54;
14'h305e:data=8'h54;
14'h305f:data=8'h54;
14'h3060:data=8'h54;
14'h3061:data=8'h54;
14'h3062:data=8'h54;
14'h3063:data=8'h54;
14'h3064:data=8'h54;
14'h3065:data=8'h54;
14'h3066:data=8'h54;
14'h3067:data=8'h54;
14'h3068:data=8'h54;
14'h3069:data=8'h54;
14'h306a:data=8'h54;
14'h306b:data=8'h54;
14'h306c:data=8'h54;
14'h306d:data=8'h54;
14'h306e:data=8'h54;
14'h306f:data=8'h54;
14'h3070:data=8'h54;
14'h3071:data=8'h54;
14'h3072:data=8'h54;
14'h3073:data=8'h50;
14'h3074:data=8'h50;
14'h3075:data=8'h50;
14'h3076:data=8'h50;
14'h3077:data=8'h50;
14'h3078:data=8'h40;
14'h3079:data=8'h40;
14'h307a:data=8'h40;
14'h307b:data=8'h40;
14'h307c:data=8'h40;
14'h307d:data=8'h00;
14'h307e:data=8'h00;
14'h307f:data=8'h00;
14'h3800:data=8'h00;
14'h3801:data=8'h00;
14'h3802:data=8'h00;
14'h3803:data=8'h00;
14'h3804:data=8'h00;
14'h3805:data=8'h00;
14'h3806:data=8'h00;
14'h3807:data=8'h00;
14'h3808:data=8'h00;
14'h3809:data=8'h00;
14'h380a:data=8'h00;
14'h380b:data=8'h00;
14'h380c:data=8'h00;
14'h380d:data=8'h00;
14'h380e:data=8'h00;
14'h380f:data=8'h00;
14'h3810:data=8'h00;
14'h3811:data=8'h00;
14'h3812:data=8'h00;
14'h3813:data=8'h00;
14'h3814:data=8'h00;
14'h3815:data=8'h00;
14'h3816:data=8'h00;
14'h3817:data=8'h00;
14'h3818:data=8'h00;
14'h3819:data=8'h00;
14'h381a:data=8'h00;
14'h381b:data=8'h00;
14'h381c:data=8'h00;
14'h381d:data=8'h00;
14'h381e:data=8'h00;
14'h381f:data=8'h00;
14'h3820:data=8'h00;
14'h3821:data=8'h00;
14'h3822:data=8'h00;
14'h3823:data=8'h00;
14'h3824:data=8'h00;
14'h3825:data=8'h00;
14'h3826:data=8'h00;
14'h3827:data=8'h00;
14'h3828:data=8'h00;
14'h3829:data=8'h00;
14'h382a:data=8'h00;
14'h382b:data=8'h00;
14'h382c:data=8'h00;
14'h382d:data=8'h00;
14'h382e:data=8'h00;
14'h382f:data=8'h00;
14'h3830:data=8'h00;
14'h3831:data=8'h00;
14'h3832:data=8'h00;
14'h3833:data=8'h00;
14'h3834:data=8'h00;
14'h3835:data=8'h00;
14'h3836:data=8'h00;
14'h3837:data=8'h00;
14'h3838:data=8'h00;
14'h3839:data=8'h00;
14'h383a:data=8'h00;
14'h383b:data=8'h00;
14'h383c:data=8'h00;
14'h383d:data=8'h00;
14'h383e:data=8'h00;
14'h383f:data=8'h00;
14'h3840:data=8'h00;
14'h3841:data=8'h00;
14'h3842:data=8'h00;
14'h3843:data=8'h00;
14'h3844:data=8'h00;
14'h3845:data=8'h00;
14'h3846:data=8'h00;
14'h3847:data=8'h00;
14'h3848:data=8'h00;
14'h3849:data=8'h00;
14'h384a:data=8'h00;
14'h384b:data=8'h00;
14'h384c:data=8'h00;
14'h384d:data=8'h00;
14'h384e:data=8'h00;
14'h384f:data=8'h00;
14'h3850:data=8'h00;
14'h3851:data=8'h00;
14'h3852:data=8'h00;
14'h3853:data=8'h00;
14'h3854:data=8'h00;
14'h3855:data=8'h00;
14'h3856:data=8'h00;
14'h3857:data=8'h00;
14'h3858:data=8'h00;
14'h3859:data=8'h00;
14'h385a:data=8'h00;
14'h385b:data=8'h00;
14'h385c:data=8'h00;
14'h385d:data=8'h00;
14'h385e:data=8'h00;
14'h385f:data=8'h00;
14'h3860:data=8'h00;
14'h3861:data=8'h00;
14'h3862:data=8'h00;
14'h3863:data=8'h00;
14'h3864:data=8'h00;
14'h3865:data=8'h00;
14'h3866:data=8'h00;
14'h3867:data=8'h00;
14'h3868:data=8'h00;
14'h3869:data=8'h00;
14'h386a:data=8'h00;
14'h386b:data=8'h00;
14'h386c:data=8'h00;
14'h386d:data=8'h00;
14'h386e:data=8'h00;
14'h386f:data=8'h00;
14'h3870:data=8'h00;
14'h3871:data=8'h00;
14'h3872:data=8'h00;
14'h3873:data=8'h00;
14'h3874:data=8'h00;
14'h3875:data=8'h00;
14'h3876:data=8'h00;
14'h3877:data=8'h00;
14'h3878:data=8'h00;
14'h3879:data=8'h00;
14'h387a:data=8'h00;
14'h387b:data=8'h00;
14'h387c:data=8'h00;
14'h387d:data=8'h00;
14'h387e:data=8'h00;
14'h387f:data=8'h00;
/////////////////////////////////////////////////////////////////////////PIC2 Dire
14'h0100:data=8'h00;
14'h0101:data=8'h00;
14'h0102:data=8'h00;
14'h0103:data=8'h00;
14'h0104:data=8'h00;
14'h0105:data=8'h00;
14'h0106:data=8'h00;
14'h0107:data=8'h00;
14'h0108:data=8'h00;
14'h0109:data=8'h00;
14'h010a:data=8'h00;
14'h010b:data=8'h00;
14'h010c:data=8'h00;
14'h010d:data=8'h00;
14'h010e:data=8'h00;
14'h010f:data=8'h00;
14'h0110:data=8'h00;
14'h0111:data=8'h00;
14'h0112:data=8'h00;
14'h0113:data=8'h00;
14'h0114:data=8'h00;
14'h0115:data=8'h00;
14'h0116:data=8'h00;
14'h0117:data=8'h00;
14'h0118:data=8'h00;
14'h0119:data=8'h00;
14'h011a:data=8'h00;
14'h011b:data=8'h00;
14'h011c:data=8'h00;
14'h011d:data=8'h00;
14'h011e:data=8'h00;
14'h011f:data=8'h00;
14'h0120:data=8'h00;
14'h0121:data=8'h00;
14'h0122:data=8'h00;
14'h0123:data=8'h00;
14'h0124:data=8'h00;
14'h0125:data=8'h00;
14'h0126:data=8'h00;
14'h0127:data=8'h00;
14'h0128:data=8'h00;
14'h0129:data=8'h00;
14'h012a:data=8'h00;
14'h012b:data=8'h00;
14'h012c:data=8'h00;
14'h012d:data=8'h00;
14'h012e:data=8'h00;
14'h012f:data=8'h00;
14'h0130:data=8'h00;
14'h0131:data=8'h00;
14'h0132:data=8'h00;
14'h0133:data=8'h00;
14'h0134:data=8'h00;
14'h0135:data=8'h00;
14'h0136:data=8'h00;
14'h0137:data=8'h00;
14'h0138:data=8'h00;
14'h0139:data=8'h00;
14'h013a:data=8'h00;
14'h013b:data=8'h00;
14'h013c:data=8'h00;
14'h013d:data=8'h00;
14'h013e:data=8'h00;
14'h013f:data=8'h00;
14'h0140:data=8'h00;
14'h0141:data=8'h00;
14'h0142:data=8'h00;
14'h0143:data=8'h00;
14'h0144:data=8'h00;
14'h0145:data=8'h00;
14'h0146:data=8'h00;
14'h0147:data=8'h00;
14'h0148:data=8'h00;
14'h0149:data=8'h00;
14'h014a:data=8'h00;
14'h014b:data=8'h00;
14'h014c:data=8'h00;
14'h014d:data=8'h00;
14'h014e:data=8'h00;
14'h014f:data=8'h00;
14'h0150:data=8'h00;
14'h0151:data=8'h00;
14'h0152:data=8'h00;
14'h0153:data=8'h00;
14'h0154:data=8'h00;
14'h0155:data=8'h00;
14'h0156:data=8'h00;
14'h0157:data=8'h00;
14'h0158:data=8'h00;
14'h0159:data=8'h00;
14'h015a:data=8'h00;
14'h015b:data=8'h00;
14'h015c:data=8'h00;
14'h015d:data=8'h00;
14'h015e:data=8'h00;
14'h015f:data=8'h00;
14'h0160:data=8'h00;
14'h0161:data=8'h00;
14'h0162:data=8'h00;
14'h0163:data=8'h00;
14'h0164:data=8'h00;
14'h0165:data=8'h00;
14'h0166:data=8'h00;
14'h0167:data=8'h00;
14'h0168:data=8'h00;
14'h0169:data=8'h00;
14'h016a:data=8'h00;
14'h016b:data=8'h00;
14'h016c:data=8'h00;
14'h016d:data=8'h00;
14'h016e:data=8'h00;
14'h016f:data=8'h00;
14'h0170:data=8'h00;
14'h0171:data=8'h00;
14'h0172:data=8'h00;
14'h0173:data=8'h00;
14'h0174:data=8'h00;
14'h0175:data=8'h00;
14'h0176:data=8'h00;
14'h0177:data=8'h00;
14'h0178:data=8'h00;
14'h0179:data=8'h00;
14'h017a:data=8'h00;
14'h017b:data=8'h00;
14'h017c:data=8'h00;
14'h017d:data=8'h00;
14'h017e:data=8'h00;
14'h017f:data=8'h00;
14'h0900:data=8'h00;
14'h0901:data=8'h00;
14'h0902:data=8'h00;
14'h0903:data=8'h00;
14'h0904:data=8'h00;
14'h0905:data=8'h00;
14'h0906:data=8'h00;
14'h0907:data=8'h00;
14'h0908:data=8'h00;
14'h0909:data=8'h00;
14'h090a:data=8'h00;
14'h090b:data=8'h00;
14'h090c:data=8'h00;
14'h090d:data=8'h00;
14'h090e:data=8'h00;
14'h090f:data=8'h00;
14'h0910:data=8'h00;
14'h0911:data=8'h00;
14'h0912:data=8'h00;
14'h0913:data=8'h00;
14'h0914:data=8'h00;
14'h0915:data=8'h00;
14'h0916:data=8'h00;
14'h0917:data=8'h00;
14'h0918:data=8'h00;
14'h0919:data=8'h00;
14'h091a:data=8'h00;
14'h091b:data=8'h00;
14'h091c:data=8'h00;
14'h091d:data=8'h00;
14'h091e:data=8'h00;
14'h091f:data=8'h00;
14'h0920:data=8'h00;
14'h0921:data=8'h00;
14'h0922:data=8'h00;
14'h0923:data=8'h00;
14'h0924:data=8'h00;
14'h0925:data=8'h00;
14'h0926:data=8'h00;
14'h0927:data=8'h00;
14'h0928:data=8'h00;
14'h0929:data=8'h00;
14'h092a:data=8'h00;
14'h092b:data=8'h00;
14'h092c:data=8'h00;
14'h092d:data=8'h00;
14'h092e:data=8'h00;
14'h092f:data=8'h00;
14'h0930:data=8'h00;
14'h0931:data=8'h00;
14'h0932:data=8'h00;
14'h0933:data=8'h00;
14'h0934:data=8'h00;
14'h0935:data=8'h00;
14'h0936:data=8'h00;
14'h0937:data=8'h00;
14'h0938:data=8'h00;
14'h0939:data=8'h80;
14'h093a:data=8'h80;
14'h093b:data=8'h80;
14'h093c:data=8'h80;
14'h093d:data=8'h80;
14'h093e:data=8'h80;
14'h093f:data=8'h80;
14'h0940:data=8'h00;
14'h0941:data=8'h00;
14'h0942:data=8'h00;
14'h0943:data=8'h00;
14'h0944:data=8'h00;
14'h0945:data=8'h00;
14'h0946:data=8'h00;
14'h0947:data=8'h00;
14'h0948:data=8'h00;
14'h0949:data=8'h00;
14'h094a:data=8'h00;
14'h094b:data=8'h00;
14'h094c:data=8'h00;
14'h094d:data=8'h00;
14'h094e:data=8'h00;
14'h094f:data=8'h00;
14'h0950:data=8'h00;
14'h0951:data=8'h00;
14'h0952:data=8'h00;
14'h0953:data=8'h00;
14'h0954:data=8'h00;
14'h0955:data=8'h00;
14'h0956:data=8'h00;
14'h0957:data=8'h00;
14'h0958:data=8'h00;
14'h0959:data=8'h00;
14'h095a:data=8'h00;
14'h095b:data=8'h00;
14'h095c:data=8'h00;
14'h095d:data=8'h00;
14'h095e:data=8'h00;
14'h095f:data=8'h00;
14'h0960:data=8'h00;
14'h0961:data=8'h00;
14'h0962:data=8'h00;
14'h0963:data=8'h00;
14'h0964:data=8'h00;
14'h0965:data=8'h00;
14'h0966:data=8'h00;
14'h0967:data=8'h00;
14'h0968:data=8'h00;
14'h0969:data=8'h00;
14'h096a:data=8'h00;
14'h096b:data=8'h00;
14'h096c:data=8'h00;
14'h096d:data=8'h00;
14'h096e:data=8'h00;
14'h096f:data=8'h00;
14'h0970:data=8'h00;
14'h0971:data=8'h00;
14'h0972:data=8'h00;
14'h0973:data=8'h00;
14'h0974:data=8'h00;
14'h0975:data=8'h00;
14'h0976:data=8'h00;
14'h0977:data=8'h00;
14'h0978:data=8'h00;
14'h0979:data=8'h00;
14'h097a:data=8'h00;
14'h097b:data=8'h00;
14'h097c:data=8'h00;
14'h097d:data=8'h00;
14'h097e:data=8'h00;
14'h097f:data=8'h00;
14'h1100:data=8'h00;
14'h1101:data=8'h00;
14'h1102:data=8'h00;
14'h1103:data=8'h00;
14'h1104:data=8'h00;
14'h1105:data=8'h00;
14'h1106:data=8'h00;
14'h1107:data=8'h00;
14'h1108:data=8'h00;
14'h1109:data=8'h00;
14'h110a:data=8'h00;
14'h110b:data=8'h00;
14'h110c:data=8'h00;
14'h110d:data=8'h00;
14'h110e:data=8'h00;
14'h110f:data=8'h00;
14'h1110:data=8'h00;
14'h1111:data=8'h00;
14'h1112:data=8'h00;
14'h1113:data=8'h00;
14'h1114:data=8'h00;
14'h1115:data=8'h00;
14'h1116:data=8'h00;
14'h1117:data=8'h00;
14'h1118:data=8'h00;
14'h1119:data=8'hF8;
14'h111a:data=8'hFE;
14'h111b:data=8'hFE;
14'h111c:data=8'hFE;
14'h111d:data=8'hFE;
14'h111e:data=8'hFE;
14'h111f:data=8'hFE;
14'h1120:data=8'hFE;
14'h1121:data=8'hFE;
14'h1122:data=8'hFE;
14'h1123:data=8'hFE;
14'h1124:data=8'hFE;
14'h1125:data=8'hFE;
14'h1126:data=8'hFE;
14'h1127:data=8'hFE;
14'h1128:data=8'hFE;
14'h1129:data=8'hFE;
14'h112a:data=8'hFE;
14'h112b:data=8'hFE;
14'h112c:data=8'hFC;
14'h112d:data=8'hFC;
14'h112e:data=8'hF8;
14'h112f:data=8'hF0;
14'h1130:data=8'hE0;
14'h1131:data=8'hC0;
14'h1132:data=8'h00;
14'h1133:data=8'h00;
14'h1134:data=8'h00;
14'h1135:data=8'h00;
14'h1136:data=8'h00;
14'h1137:data=8'h00;
14'h1138:data=8'h3F;
14'h1139:data=8'h7F;
14'h113a:data=8'hFF;
14'h113b:data=8'hFF;
14'h113c:data=8'hFF;
14'h113d:data=8'hFF;
14'h113e:data=8'hFF;
14'h113f:data=8'h7F;
14'h1140:data=8'h3F;
14'h1141:data=8'h00;
14'h1142:data=8'h00;
14'h1143:data=8'h00;
14'h1144:data=8'h00;
14'h1145:data=8'h00;
14'h1146:data=8'h00;
14'h1147:data=8'h00;
14'h1148:data=8'h00;
14'h1149:data=8'h00;
14'h114a:data=8'h00;
14'h114b:data=8'h00;
14'h114c:data=8'h00;
14'h114d:data=8'h00;
14'h114e:data=8'h00;
14'h114f:data=8'h00;
14'h1150:data=8'h00;
14'h1151:data=8'h00;
14'h1152:data=8'h00;
14'h1153:data=8'h00;
14'h1154:data=8'h00;
14'h1155:data=8'h00;
14'h1156:data=8'h00;
14'h1157:data=8'h00;
14'h1158:data=8'h00;
14'h1159:data=8'h00;
14'h115a:data=8'h00;
14'h115b:data=8'h00;
14'h115c:data=8'h00;
14'h115d:data=8'h00;
14'h115e:data=8'h00;
14'h115f:data=8'h00;
14'h1160:data=8'h00;
14'h1161:data=8'h00;
14'h1162:data=8'h00;
14'h1163:data=8'h00;
14'h1164:data=8'h00;
14'h1165:data=8'h00;
14'h1166:data=8'h00;
14'h1167:data=8'h00;
14'h1168:data=8'h00;
14'h1169:data=8'h00;
14'h116a:data=8'h00;
14'h116b:data=8'h00;
14'h116c:data=8'h00;
14'h116d:data=8'h00;
14'h116e:data=8'h00;
14'h116f:data=8'h00;
14'h1170:data=8'h00;
14'h1171:data=8'h00;
14'h1172:data=8'h00;
14'h1173:data=8'h00;
14'h1174:data=8'h00;
14'h1175:data=8'h00;
14'h1176:data=8'h00;
14'h1177:data=8'h00;
14'h1178:data=8'h00;
14'h1179:data=8'h00;
14'h117a:data=8'h00;
14'h117b:data=8'h00;
14'h117c:data=8'h00;
14'h117d:data=8'h00;
14'h117e:data=8'h00;
14'h117f:data=8'h00;
14'h1900:data=8'h00;
14'h1901:data=8'h00;
14'h1902:data=8'h00;
14'h1903:data=8'h00;
14'h1904:data=8'h00;
14'h1905:data=8'h00;
14'h1906:data=8'h00;
14'h1907:data=8'h00;
14'h1908:data=8'h00;
14'h1909:data=8'h00;
14'h190a:data=8'h00;
14'h190b:data=8'h00;
14'h190c:data=8'h00;
14'h190d:data=8'h00;
14'h190e:data=8'h00;
14'h190f:data=8'h00;
14'h1910:data=8'h00;
14'h1911:data=8'h00;
14'h1912:data=8'h00;
14'h1913:data=8'h00;
14'h1914:data=8'h00;
14'h1915:data=8'h00;
14'h1916:data=8'h00;
14'h1917:data=8'hE0;
14'h1918:data=8'hFF;
14'h1919:data=8'hFF;
14'h191a:data=8'hFF;
14'h191b:data=8'hFF;
14'h191c:data=8'hFF;
14'h191d:data=8'hFF;
14'h191e:data=8'hFF;
14'h191f:data=8'hFF;
14'h1920:data=8'h07;
14'h1921:data=8'h00;
14'h1922:data=8'h00;
14'h1923:data=8'h00;
14'h1924:data=8'h00;
14'h1925:data=8'h00;
14'h1926:data=8'h01;
14'h1927:data=8'h01;
14'h1928:data=8'h03;
14'h1929:data=8'h03;
14'h192a:data=8'hFF;
14'h192b:data=8'hFF;
14'h192c:data=8'hFF;
14'h192d:data=8'hFF;
14'h192e:data=8'hFF;
14'h192f:data=8'hFF;
14'h1930:data=8'hFF;
14'h1931:data=8'hFF;
14'h1932:data=8'hFE;
14'h1933:data=8'h00;
14'h1934:data=8'h00;
14'h1935:data=8'h80;
14'h1936:data=8'hF8;
14'h1937:data=8'hFE;
14'h1938:data=8'hFE;
14'h1939:data=8'hFE;
14'h193a:data=8'hFE;
14'h193b:data=8'hFE;
14'h193c:data=8'hFE;
14'h193d:data=8'hFE;
14'h193e:data=8'h7E;
14'h193f:data=8'h00;
14'h1940:data=8'h00;
14'h1941:data=8'h00;
14'h1942:data=8'h00;
14'h1943:data=8'hE0;
14'h1944:data=8'hFE;
14'h1945:data=8'hFE;
14'h1946:data=8'hFE;
14'h1947:data=8'hFE;
14'h1948:data=8'hFE;
14'h1949:data=8'hFE;
14'h194a:data=8'hFE;
14'h194b:data=8'hFE;
14'h194c:data=8'hFC;
14'h194d:data=8'hFE;
14'h194e:data=8'hFE;
14'h194f:data=8'hFE;
14'h1950:data=8'hFE;
14'h1951:data=8'hFE;
14'h1952:data=8'hFE;
14'h1953:data=8'h9E;
14'h1954:data=8'hE0;
14'h1955:data=8'hF0;
14'h1956:data=8'hF8;
14'h1957:data=8'hF8;
14'h1958:data=8'hFC;
14'h1959:data=8'hFC;
14'h195a:data=8'hFE;
14'h195b:data=8'hFE;
14'h195c:data=8'hFE;
14'h195d:data=8'hFE;
14'h195e:data=8'h7E;
14'h195f:data=8'hFE;
14'h1960:data=8'hFE;
14'h1961:data=8'hFE;
14'h1962:data=8'hFE;
14'h1963:data=8'hFE;
14'h1964:data=8'hFE;
14'h1965:data=8'hFC;
14'h1966:data=8'hF8;
14'h1967:data=8'hE0;
14'h1968:data=8'h00;
14'h1969:data=8'h00;
14'h196a:data=8'h00;
14'h196b:data=8'h00;
14'h196c:data=8'h00;
14'h196d:data=8'h00;
14'h196e:data=8'h00;
14'h196f:data=8'h00;
14'h1970:data=8'h00;
14'h1971:data=8'h00;
14'h1972:data=8'h00;
14'h1973:data=8'h00;
14'h1974:data=8'h00;
14'h1975:data=8'h00;
14'h1976:data=8'h00;
14'h1977:data=8'h00;
14'h1978:data=8'h00;
14'h1979:data=8'h00;
14'h197a:data=8'h00;
14'h197b:data=8'h00;
14'h197c:data=8'h00;
14'h197d:data=8'h00;
14'h197e:data=8'h00;
14'h197f:data=8'h00;
14'h2100:data=8'h00;
14'h2101:data=8'h00;
14'h2102:data=8'h00;
14'h2103:data=8'h00;
14'h2104:data=8'h00;
14'h2105:data=8'h00;
14'h2106:data=8'h00;
14'h2107:data=8'h00;
14'h2108:data=8'h00;
14'h2109:data=8'h00;
14'h210a:data=8'h00;
14'h210b:data=8'h00;
14'h210c:data=8'h00;
14'h210d:data=8'h00;
14'h210e:data=8'h00;
14'h210f:data=8'h00;
14'h2110:data=8'h00;
14'h2111:data=8'h00;
14'h2112:data=8'h00;
14'h2113:data=8'h00;
14'h2114:data=8'h00;
14'h2115:data=8'hC0;
14'h2116:data=8'hFE;
14'h2117:data=8'hFF;
14'h2118:data=8'hFF;
14'h2119:data=8'hFF;
14'h211a:data=8'hFF;
14'h211b:data=8'hFF;
14'h211c:data=8'hFF;
14'h211d:data=8'hFF;
14'h211e:data=8'h1F;
14'h211f:data=8'h00;
14'h2120:data=8'h00;
14'h2121:data=8'h00;
14'h2122:data=8'h00;
14'h2123:data=8'h00;
14'h2124:data=8'h00;
14'h2125:data=8'h00;
14'h2126:data=8'h80;
14'h2127:data=8'hC0;
14'h2128:data=8'hE0;
14'h2129:data=8'hF8;
14'h212a:data=8'hFF;
14'h212b:data=8'hFF;
14'h212c:data=8'hFF;
14'h212d:data=8'hFF;
14'h212e:data=8'hFF;
14'h212f:data=8'hFF;
14'h2130:data=8'hFF;
14'h2131:data=8'h7F;
14'h2132:data=8'h0F;
14'h2133:data=8'h00;
14'h2134:data=8'hF0;
14'h2135:data=8'hFF;
14'h2136:data=8'hFF;
14'h2137:data=8'hFF;
14'h2138:data=8'hFF;
14'h2139:data=8'hFF;
14'h213a:data=8'hFF;
14'h213b:data=8'hFF;
14'h213c:data=8'hFF;
14'h213d:data=8'h07;
14'h213e:data=8'h00;
14'h213f:data=8'h00;
14'h2140:data=8'h00;
14'h2141:data=8'h80;
14'h2142:data=8'hFC;
14'h2143:data=8'hFF;
14'h2144:data=8'hFF;
14'h2145:data=8'hFF;
14'h2146:data=8'hFF;
14'h2147:data=8'hFF;
14'h2148:data=8'hFF;
14'h2149:data=8'hFF;
14'h214a:data=8'h3F;
14'h214b:data=8'h0F;
14'h214c:data=8'h07;
14'h214d:data=8'h03;
14'h214e:data=8'h01;
14'h214f:data=8'h01;
14'h2150:data=8'h01;
14'h2151:data=8'h03;
14'h2152:data=8'hFF;
14'h2153:data=8'hFF;
14'h2154:data=8'hFF;
14'h2155:data=8'hFF;
14'h2156:data=8'hFF;
14'h2157:data=8'hFF;
14'h2158:data=8'hFF;
14'h2159:data=8'hFF;
14'h215a:data=8'hFF;
14'h215b:data=8'hFF;
14'h215c:data=8'hFE;
14'h215d:data=8'hFE;
14'h215e:data=8'hFF;
14'h215f:data=8'hFF;
14'h2160:data=8'h7F;
14'h2161:data=8'h7F;
14'h2162:data=8'h7F;
14'h2163:data=8'hFF;
14'h2164:data=8'hBF;
14'h2165:data=8'h1F;
14'h2166:data=8'h0F;
14'h2167:data=8'h03;
14'h2168:data=8'h00;
14'h2169:data=8'h00;
14'h216a:data=8'h00;
14'h216b:data=8'h00;
14'h216c:data=8'h00;
14'h216d:data=8'h00;
14'h216e:data=8'h00;
14'h216f:data=8'h00;
14'h2170:data=8'h00;
14'h2171:data=8'h00;
14'h2172:data=8'h00;
14'h2173:data=8'h00;
14'h2174:data=8'h00;
14'h2175:data=8'h00;
14'h2176:data=8'h00;
14'h2177:data=8'h00;
14'h2178:data=8'h00;
14'h2179:data=8'h00;
14'h217a:data=8'h00;
14'h217b:data=8'h00;
14'h217c:data=8'h00;
14'h217d:data=8'h00;
14'h217e:data=8'h00;
14'h217f:data=8'h00;
14'h2900:data=8'h00;
14'h2901:data=8'h00;
14'h2902:data=8'h00;
14'h2903:data=8'h00;
14'h2904:data=8'h00;
14'h2905:data=8'h00;
14'h2906:data=8'h00;
14'h2907:data=8'h00;
14'h2908:data=8'h00;
14'h2909:data=8'h00;
14'h290a:data=8'h00;
14'h290b:data=8'h00;
14'h290c:data=8'h00;
14'h290d:data=8'h00;
14'h290e:data=8'h00;
14'h290f:data=8'h00;
14'h2910:data=8'h00;
14'h2911:data=8'h00;
14'h2912:data=8'h00;
14'h2913:data=8'h00;
14'h2914:data=8'h00;
14'h2915:data=8'hFF;
14'h2916:data=8'hFF;
14'h2917:data=8'hFF;
14'h2918:data=8'hFF;
14'h2919:data=8'hFF;
14'h291a:data=8'hFF;
14'h291b:data=8'hFF;
14'h291c:data=8'hFF;
14'h291d:data=8'hFF;
14'h291e:data=8'hFC;
14'h291f:data=8'hFC;
14'h2920:data=8'hFC;
14'h2921:data=8'hFC;
14'h2922:data=8'hFE;
14'h2923:data=8'hFE;
14'h2924:data=8'hFF;
14'h2925:data=8'hFF;
14'h2926:data=8'hFF;
14'h2927:data=8'hFF;
14'h2928:data=8'h7F;
14'h2929:data=8'h7F;
14'h292a:data=8'h3F;
14'h292b:data=8'h3F;
14'h292c:data=8'h1F;
14'h292d:data=8'h0F;
14'h292e:data=8'h07;
14'h292f:data=8'h03;
14'h2930:data=8'h01;
14'h2931:data=8'h00;
14'h2932:data=8'h00;
14'h2933:data=8'h00;
14'h2934:data=8'h1F;
14'h2935:data=8'h7F;
14'h2936:data=8'h7F;
14'h2937:data=8'hFF;
14'h2938:data=8'hFF;
14'h2939:data=8'hFF;
14'h293a:data=8'hFF;
14'h293b:data=8'hFF;
14'h293c:data=8'hFE;
14'h293d:data=8'hFE;
14'h293e:data=8'hFE;
14'h293f:data=8'h1E;
14'h2940:data=8'hF0;
14'h2941:data=8'hFF;
14'h2942:data=8'hFF;
14'h2943:data=8'hFF;
14'h2944:data=8'hFF;
14'h2945:data=8'hFF;
14'h2946:data=8'hFF;
14'h2947:data=8'hFF;
14'h2948:data=8'h7F;
14'h2949:data=8'h03;
14'h294a:data=8'h00;
14'h294b:data=8'h00;
14'h294c:data=8'h00;
14'h294d:data=8'h00;
14'h294e:data=8'h00;
14'h294f:data=8'h00;
14'h2950:data=8'h00;
14'h2951:data=8'h00;
14'h2952:data=8'h07;
14'h2953:data=8'h1F;
14'h2954:data=8'h3F;
14'h2955:data=8'h7F;
14'h2956:data=8'h7F;
14'h2957:data=8'hFF;
14'h2958:data=8'hFF;
14'h2959:data=8'hFF;
14'h295a:data=8'hFF;
14'h295b:data=8'hFE;
14'h295c:data=8'hFE;
14'h295d:data=8'hFC;
14'h295e:data=8'hFE;
14'h295f:data=8'hFE;
14'h2960:data=8'hFE;
14'h2961:data=8'hFF;
14'h2962:data=8'h7F;
14'h2963:data=8'h7F;
14'h2964:data=8'h07;
14'h2965:data=8'h00;
14'h2966:data=8'h00;
14'h2967:data=8'h00;
14'h2968:data=8'h00;
14'h2969:data=8'h00;
14'h296a:data=8'h00;
14'h296b:data=8'h00;
14'h296c:data=8'h00;
14'h296d:data=8'h00;
14'h296e:data=8'h00;
14'h296f:data=8'h00;
14'h2970:data=8'h00;
14'h2971:data=8'h00;
14'h2972:data=8'h00;
14'h2973:data=8'h00;
14'h2974:data=8'h00;
14'h2975:data=8'h00;
14'h2976:data=8'h00;
14'h2977:data=8'h00;
14'h2978:data=8'h00;
14'h2979:data=8'h00;
14'h297a:data=8'h00;
14'h297b:data=8'h00;
14'h297c:data=8'h00;
14'h297d:data=8'h00;
14'h297e:data=8'h00;
14'h297f:data=8'h00;
14'h3100:data=8'h00;
14'h3101:data=8'h00;
14'h3102:data=8'h00;
14'h3103:data=8'h00;
14'h3104:data=8'h00;
14'h3105:data=8'h00;
14'h3106:data=8'h00;
14'h3107:data=8'h00;
14'h3108:data=8'h00;
14'h3109:data=8'h00;
14'h310a:data=8'h00;
14'h310b:data=8'h00;
14'h310c:data=8'h00;
14'h310d:data=8'h00;
14'h310e:data=8'h00;
14'h310f:data=8'h00;
14'h3110:data=8'h00;
14'h3111:data=8'h00;
14'h3112:data=8'h00;
14'h3113:data=8'h00;
14'h3114:data=8'h00;
14'h3115:data=8'h00;
14'h3116:data=8'h00;
14'h3117:data=8'h00;
14'h3118:data=8'h00;
14'h3119:data=8'h00;
14'h311a:data=8'h00;
14'h311b:data=8'h00;
14'h311c:data=8'h00;
14'h311d:data=8'h00;
14'h311e:data=8'h00;
14'h311f:data=8'h00;
14'h3120:data=8'h00;
14'h3121:data=8'h00;
14'h3122:data=8'h00;
14'h3123:data=8'h00;
14'h3124:data=8'h00;
14'h3125:data=8'h00;
14'h3126:data=8'h00;
14'h3127:data=8'h00;
14'h3128:data=8'h00;
14'h3129:data=8'h00;
14'h312a:data=8'h00;
14'h312b:data=8'h00;
14'h312c:data=8'h00;
14'h312d:data=8'h00;
14'h312e:data=8'h00;
14'h312f:data=8'h00;
14'h3130:data=8'h00;
14'h3131:data=8'h00;
14'h3132:data=8'h00;
14'h3133:data=8'h00;
14'h3134:data=8'h00;
14'h3135:data=8'h00;
14'h3136:data=8'h00;
14'h3137:data=8'h00;
14'h3138:data=8'h00;
14'h3139:data=8'h00;
14'h313a:data=8'h00;
14'h313b:data=8'h00;
14'h313c:data=8'h00;
14'h313d:data=8'h00;
14'h313e:data=8'h00;
14'h313f:data=8'h00;
14'h3140:data=8'h00;
14'h3141:data=8'h00;
14'h3142:data=8'h00;
14'h3143:data=8'h00;
14'h3144:data=8'h00;
14'h3145:data=8'h00;
14'h3146:data=8'h00;
14'h3147:data=8'h00;
14'h3148:data=8'h00;
14'h3149:data=8'h00;
14'h314a:data=8'h00;
14'h314b:data=8'h00;
14'h314c:data=8'h00;
14'h314d:data=8'h00;
14'h314e:data=8'h00;
14'h314f:data=8'h00;
14'h3150:data=8'h00;
14'h3151:data=8'h00;
14'h3152:data=8'h00;
14'h3153:data=8'h00;
14'h3154:data=8'h00;
14'h3155:data=8'h00;
14'h3156:data=8'h00;
14'h3157:data=8'h00;
14'h3158:data=8'h00;
14'h3159:data=8'h00;
14'h315a:data=8'h00;
14'h315b:data=8'h00;
14'h315c:data=8'h00;
14'h315d:data=8'h00;
14'h315e:data=8'h00;
14'h315f:data=8'h00;
14'h3160:data=8'h00;
14'h3161:data=8'h00;
14'h3162:data=8'h00;
14'h3163:data=8'h00;
14'h3164:data=8'h00;
14'h3165:data=8'h00;
14'h3166:data=8'h00;
14'h3167:data=8'h00;
14'h3168:data=8'h00;
14'h3169:data=8'h00;
14'h316a:data=8'h00;
14'h316b:data=8'h00;
14'h316c:data=8'h00;
14'h316d:data=8'h00;
14'h316e:data=8'h00;
14'h316f:data=8'h00;
14'h3170:data=8'h00;
14'h3171:data=8'h00;
14'h3172:data=8'h00;
14'h3173:data=8'h00;
14'h3174:data=8'h00;
14'h3175:data=8'h00;
14'h3176:data=8'h00;
14'h3177:data=8'h00;
14'h3178:data=8'h00;
14'h3179:data=8'h00;
14'h317a:data=8'h00;
14'h317b:data=8'h00;
14'h317c:data=8'h00;
14'h317d:data=8'h00;
14'h317e:data=8'h00;
14'h317f:data=8'h00;
14'h3900:data=8'h00;
14'h3901:data=8'h00;
14'h3902:data=8'h00;
14'h3903:data=8'h00;
14'h3904:data=8'h00;
14'h3905:data=8'h00;
14'h3906:data=8'h00;
14'h3907:data=8'h00;
14'h3908:data=8'h00;
14'h3909:data=8'h00;
14'h390a:data=8'h00;
14'h390b:data=8'h00;
14'h390c:data=8'h00;
14'h390d:data=8'h00;
14'h390e:data=8'h00;
14'h390f:data=8'h00;
14'h3910:data=8'h00;
14'h3911:data=8'h00;
14'h3912:data=8'h00;
14'h3913:data=8'h00;
14'h3914:data=8'h00;
14'h3915:data=8'h00;
14'h3916:data=8'h00;
14'h3917:data=8'h00;
14'h3918:data=8'h00;
14'h3919:data=8'h00;
14'h391a:data=8'h00;
14'h391b:data=8'h00;
14'h391c:data=8'h00;
14'h391d:data=8'h00;
14'h391e:data=8'h00;
14'h391f:data=8'h00;
14'h3920:data=8'h00;
14'h3921:data=8'h00;
14'h3922:data=8'h00;
14'h3923:data=8'h00;
14'h3924:data=8'h00;
14'h3925:data=8'h00;
14'h3926:data=8'h00;
14'h3927:data=8'h00;
14'h3928:data=8'h00;
14'h3929:data=8'h00;
14'h392a:data=8'h00;
14'h392b:data=8'h00;
14'h392c:data=8'h00;
14'h392d:data=8'h00;
14'h392e:data=8'h00;
14'h392f:data=8'h00;
14'h3930:data=8'h00;
14'h3931:data=8'h00;
14'h3932:data=8'h00;
14'h3933:data=8'h00;
14'h3934:data=8'h00;
14'h3935:data=8'h00;
14'h3936:data=8'h00;
14'h3937:data=8'h00;
14'h3938:data=8'h00;
14'h3939:data=8'h00;
14'h393a:data=8'h00;
14'h393b:data=8'h00;
14'h393c:data=8'h00;
14'h393d:data=8'h00;
14'h393e:data=8'h00;
14'h393f:data=8'h00;
14'h3940:data=8'h00;
14'h3941:data=8'h00;
14'h3942:data=8'h00;
14'h3943:data=8'h00;
14'h3944:data=8'h00;
14'h3945:data=8'h00;
14'h3946:data=8'h00;
14'h3947:data=8'h00;
14'h3948:data=8'h00;
14'h3949:data=8'h00;
14'h394a:data=8'h00;
14'h394b:data=8'h00;
14'h394c:data=8'h00;
14'h394d:data=8'h00;
14'h394e:data=8'h00;
14'h394f:data=8'h00;
14'h3950:data=8'h00;
14'h3951:data=8'h00;
14'h3952:data=8'h00;
14'h3953:data=8'h00;
14'h3954:data=8'h00;
14'h3955:data=8'h00;
14'h3956:data=8'h00;
14'h3957:data=8'h00;
14'h3958:data=8'h00;
14'h3959:data=8'h00;
14'h395a:data=8'h00;
14'h395b:data=8'h00;
14'h395c:data=8'h00;
14'h395d:data=8'h00;
14'h395e:data=8'h00;
14'h395f:data=8'h00;
14'h3960:data=8'h00;
14'h3961:data=8'h00;
14'h3962:data=8'h00;
14'h3963:data=8'h00;
14'h3964:data=8'h00;
14'h3965:data=8'h00;
14'h3966:data=8'h00;
14'h3967:data=8'h00;
14'h3968:data=8'h00;
14'h3969:data=8'h00;
14'h396a:data=8'h00;
14'h396b:data=8'h00;
14'h396c:data=8'h00;
14'h396d:data=8'h00;
14'h396e:data=8'h00;
14'h396f:data=8'h00;
14'h3970:data=8'h00;
14'h3971:data=8'h00;
14'h3972:data=8'h00;
14'h3973:data=8'h00;
14'h3974:data=8'h00;
14'h3975:data=8'h00;
14'h3976:data=8'h00;
14'h3977:data=8'h00;
14'h3978:data=8'h00;
14'h3979:data=8'h00;
14'h397a:data=8'h00;
14'h397b:data=8'h00;
14'h397c:data=8'h00;
14'h397d:data=8'h00;
14'h397e:data=8'h00;
14'h397f:data=8'h00;
//////////////////////////////////////////////////////////////////////PIC3 Locate
14'h0200:data=8'h00;
14'h0201:data=8'h00;
14'h0202:data=8'h00;
14'h0203:data=8'h00;
14'h0204:data=8'h00;
14'h0205:data=8'h00;
14'h0206:data=8'h00;
14'h0207:data=8'h00;
14'h0208:data=8'h00;
14'h0209:data=8'h00;
14'h020a:data=8'h00;
14'h020b:data=8'h00;
14'h020c:data=8'h00;
14'h020d:data=8'h00;
14'h020e:data=8'h00;
14'h020f:data=8'h00;
14'h0210:data=8'h00;
14'h0211:data=8'h00;
14'h0212:data=8'h00;
14'h0213:data=8'h00;
14'h0214:data=8'h00;
14'h0215:data=8'h00;
14'h0216:data=8'h00;
14'h0217:data=8'h00;
14'h0218:data=8'h00;
14'h0219:data=8'h00;
14'h021a:data=8'h00;
14'h021b:data=8'h00;
14'h021c:data=8'h00;
14'h021d:data=8'h00;
14'h021e:data=8'h00;
14'h021f:data=8'h00;
14'h0220:data=8'h00;
14'h0221:data=8'h00;
14'h0222:data=8'h00;
14'h0223:data=8'h00;
14'h0224:data=8'h00;
14'h0225:data=8'h00;
14'h0226:data=8'h00;
14'h0227:data=8'h00;
14'h0228:data=8'h00;
14'h0229:data=8'h00;
14'h022a:data=8'h00;
14'h022b:data=8'h00;
14'h022c:data=8'h00;
14'h022d:data=8'h00;
14'h022e:data=8'h00;
14'h022f:data=8'h00;
14'h0230:data=8'h00;
14'h0231:data=8'h00;
14'h0232:data=8'h00;
14'h0233:data=8'h00;
14'h0234:data=8'h00;
14'h0235:data=8'h00;
14'h0236:data=8'h00;
14'h0237:data=8'h00;
14'h0238:data=8'h00;
14'h0239:data=8'h00;
14'h023a:data=8'h00;
14'h023b:data=8'h00;
14'h023c:data=8'h00;
14'h023d:data=8'h00;
14'h023e:data=8'h00;
14'h023f:data=8'h00;
14'h0240:data=8'h00;
14'h0241:data=8'h00;
14'h0242:data=8'h00;
14'h0243:data=8'h00;
14'h0244:data=8'h00;
14'h0245:data=8'h00;
14'h0246:data=8'h00;
14'h0247:data=8'h00;
14'h0248:data=8'h00;
14'h0249:data=8'h00;
14'h024a:data=8'h00;
14'h024b:data=8'h00;
14'h024c:data=8'h00;
14'h024d:data=8'h00;
14'h024e:data=8'h00;
14'h024f:data=8'h00;
14'h0250:data=8'h00;
14'h0251:data=8'h00;
14'h0252:data=8'h00;
14'h0253:data=8'h00;
14'h0254:data=8'h00;
14'h0255:data=8'h00;
14'h0256:data=8'h00;
14'h0257:data=8'h00;
14'h0258:data=8'h00;
14'h0259:data=8'h00;
14'h025a:data=8'h00;
14'h025b:data=8'h00;
14'h025c:data=8'h00;
14'h025d:data=8'h00;
14'h025e:data=8'h00;
14'h025f:data=8'h00;
14'h0260:data=8'h00;
14'h0261:data=8'h00;
14'h0262:data=8'h00;
14'h0263:data=8'h00;
14'h0264:data=8'h00;
14'h0265:data=8'h00;
14'h0266:data=8'h00;
14'h0267:data=8'h00;
14'h0268:data=8'h00;
14'h0269:data=8'h00;
14'h026a:data=8'h00;
14'h026b:data=8'h00;
14'h026c:data=8'h00;
14'h026d:data=8'h00;
14'h026e:data=8'h00;
14'h026f:data=8'h00;
14'h0270:data=8'h00;
14'h0271:data=8'h00;
14'h0272:data=8'h00;
14'h0273:data=8'h00;
14'h0274:data=8'h00;
14'h0275:data=8'h00;
14'h0276:data=8'h00;
14'h0277:data=8'h00;
14'h0278:data=8'h00;
14'h0279:data=8'h00;
14'h027a:data=8'h00;
14'h027b:data=8'h00;
14'h027c:data=8'h00;
14'h027d:data=8'h00;
14'h027e:data=8'h00;
14'h027f:data=8'h00;
14'h0a00:data=8'h00;
14'h0a01:data=8'h00;
14'h0a02:data=8'h00;
14'h0a03:data=8'h00;
14'h0a04:data=8'h00;
14'h0a05:data=8'h00;
14'h0a06:data=8'h00;
14'h0a07:data=8'h00;
14'h0a08:data=8'h00;
14'h0a09:data=8'h00;
14'h0a0a:data=8'h00;
14'h0a0b:data=8'h00;
14'h0a0c:data=8'h00;
14'h0a0d:data=8'h00;
14'h0a0e:data=8'h00;
14'h0a0f:data=8'h00;
14'h0a10:data=8'h00;
14'h0a11:data=8'h80;
14'h0a12:data=8'hC0;
14'h0a13:data=8'hC0;
14'h0a14:data=8'hC0;
14'h0a15:data=8'hC0;
14'h0a16:data=8'hC0;
14'h0a17:data=8'hC0;
14'h0a18:data=8'hC0;
14'h0a19:data=8'h00;
14'h0a1a:data=8'h00;
14'h0a1b:data=8'h00;
14'h0a1c:data=8'h00;
14'h0a1d:data=8'h00;
14'h0a1e:data=8'h00;
14'h0a1f:data=8'h00;
14'h0a20:data=8'h00;
14'h0a21:data=8'h00;
14'h0a22:data=8'h00;
14'h0a23:data=8'h00;
14'h0a24:data=8'h00;
14'h0a25:data=8'h00;
14'h0a26:data=8'h00;
14'h0a27:data=8'h00;
14'h0a28:data=8'h00;
14'h0a29:data=8'h00;
14'h0a2a:data=8'h00;
14'h0a2b:data=8'h00;
14'h0a2c:data=8'h00;
14'h0a2d:data=8'h00;
14'h0a2e:data=8'h00;
14'h0a2f:data=8'h00;
14'h0a30:data=8'h00;
14'h0a31:data=8'h00;
14'h0a32:data=8'h00;
14'h0a33:data=8'h00;
14'h0a34:data=8'h00;
14'h0a35:data=8'h00;
14'h0a36:data=8'h00;
14'h0a37:data=8'h00;
14'h0a38:data=8'h00;
14'h0a39:data=8'h00;
14'h0a3a:data=8'h00;
14'h0a3b:data=8'h00;
14'h0a3c:data=8'h00;
14'h0a3d:data=8'h00;
14'h0a3e:data=8'h00;
14'h0a3f:data=8'h00;
14'h0a40:data=8'h00;
14'h0a41:data=8'h00;
14'h0a42:data=8'h00;
14'h0a43:data=8'h00;
14'h0a44:data=8'h00;
14'h0a45:data=8'h00;
14'h0a46:data=8'h00;
14'h0a47:data=8'h00;
14'h0a48:data=8'h00;
14'h0a49:data=8'h00;
14'h0a4a:data=8'h00;
14'h0a4b:data=8'h00;
14'h0a4c:data=8'h00;
14'h0a4d:data=8'h00;
14'h0a4e:data=8'h00;
14'h0a4f:data=8'h00;
14'h0a50:data=8'h00;
14'h0a51:data=8'h00;
14'h0a52:data=8'h00;
14'h0a53:data=8'h00;
14'h0a54:data=8'h00;
14'h0a55:data=8'h00;
14'h0a56:data=8'h00;
14'h0a57:data=8'h00;
14'h0a58:data=8'h00;
14'h0a59:data=8'h00;
14'h0a5a:data=8'h00;
14'h0a5b:data=8'h00;
14'h0a5c:data=8'h00;
14'h0a5d:data=8'h00;
14'h0a5e:data=8'h00;
14'h0a5f:data=8'h00;
14'h0a60:data=8'h00;
14'h0a61:data=8'h00;
14'h0a62:data=8'h00;
14'h0a63:data=8'h00;
14'h0a64:data=8'h00;
14'h0a65:data=8'h00;
14'h0a66:data=8'h00;
14'h0a67:data=8'h00;
14'h0a68:data=8'h00;
14'h0a69:data=8'h00;
14'h0a6a:data=8'h00;
14'h0a6b:data=8'h00;
14'h0a6c:data=8'h00;
14'h0a6d:data=8'h00;
14'h0a6e:data=8'h80;
14'h0a6f:data=8'h80;
14'h0a70:data=8'h80;
14'h0a71:data=8'h80;
14'h0a72:data=8'h80;
14'h0a73:data=8'h00;
14'h0a74:data=8'h00;
14'h0a75:data=8'h00;
14'h0a76:data=8'h00;
14'h0a77:data=8'h00;
14'h0a78:data=8'h00;
14'h0a79:data=8'h00;
14'h0a7a:data=8'h00;
14'h0a7b:data=8'h00;
14'h0a7c:data=8'h00;
14'h0a7d:data=8'h00;
14'h0a7e:data=8'h00;
14'h0a7f:data=8'h00;
14'h1200:data=8'h00;
14'h1201:data=8'h00;
14'h1202:data=8'h00;
14'h1203:data=8'h00;
14'h1204:data=8'h00;
14'h1205:data=8'h00;
14'h1206:data=8'h00;
14'h1207:data=8'h00;
14'h1208:data=8'h00;
14'h1209:data=8'h00;
14'h120a:data=8'h00;
14'h120b:data=8'h00;
14'h120c:data=8'h00;
14'h120d:data=8'h00;
14'h120e:data=8'h00;
14'h120f:data=8'hC0;
14'h1210:data=8'hFE;
14'h1211:data=8'hFF;
14'h1212:data=8'hFF;
14'h1213:data=8'hFF;
14'h1214:data=8'hFF;
14'h1215:data=8'hFF;
14'h1216:data=8'hFF;
14'h1217:data=8'hFF;
14'h1218:data=8'h0F;
14'h1219:data=8'h00;
14'h121a:data=8'h00;
14'h121b:data=8'h00;
14'h121c:data=8'h00;
14'h121d:data=8'h00;
14'h121e:data=8'h00;
14'h121f:data=8'h00;
14'h1220:data=8'h00;
14'h1221:data=8'h00;
14'h1222:data=8'h00;
14'h1223:data=8'h00;
14'h1224:data=8'h00;
14'h1225:data=8'h00;
14'h1226:data=8'h00;
14'h1227:data=8'h80;
14'h1228:data=8'h80;
14'h1229:data=8'hC0;
14'h122a:data=8'hC0;
14'h122b:data=8'hC0;
14'h122c:data=8'hC0;
14'h122d:data=8'hC0;
14'h122e:data=8'hC0;
14'h122f:data=8'hC0;
14'h1230:data=8'hC0;
14'h1231:data=8'hC0;
14'h1232:data=8'hC0;
14'h1233:data=8'h80;
14'h1234:data=8'h80;
14'h1235:data=8'h00;
14'h1236:data=8'h00;
14'h1237:data=8'h00;
14'h1238:data=8'h00;
14'h1239:data=8'h00;
14'h123a:data=8'h00;
14'h123b:data=8'h00;
14'h123c:data=8'h00;
14'h123d:data=8'h00;
14'h123e:data=8'h00;
14'h123f:data=8'h80;
14'h1240:data=8'h80;
14'h1241:data=8'hC0;
14'h1242:data=8'hC0;
14'h1243:data=8'hC0;
14'h1244:data=8'hC0;
14'h1245:data=8'hC0;
14'h1246:data=8'hC0;
14'h1247:data=8'hC0;
14'h1248:data=8'hC0;
14'h1249:data=8'hC0;
14'h124a:data=8'hC0;
14'h124b:data=8'hC0;
14'h124c:data=8'h80;
14'h124d:data=8'h00;
14'h124e:data=8'h00;
14'h124f:data=8'h00;
14'h1250:data=8'h00;
14'h1251:data=8'h00;
14'h1252:data=8'h00;
14'h1253:data=8'h80;
14'h1254:data=8'h80;
14'h1255:data=8'hC0;
14'h1256:data=8'hC0;
14'h1257:data=8'hC0;
14'h1258:data=8'hC0;
14'h1259:data=8'hC0;
14'h125a:data=8'hC0;
14'h125b:data=8'hC0;
14'h125c:data=8'hC0;
14'h125d:data=8'hC0;
14'h125e:data=8'hC0;
14'h125f:data=8'hC0;
14'h1260:data=8'hC0;
14'h1261:data=8'hC0;
14'h1262:data=8'hC0;
14'h1263:data=8'h80;
14'h1264:data=8'h80;
14'h1265:data=8'h00;
14'h1266:data=8'hC0;
14'h1267:data=8'hC0;
14'h1268:data=8'hC0;
14'h1269:data=8'hF0;
14'h126a:data=8'hFF;
14'h126b:data=8'hFF;
14'h126c:data=8'hFF;
14'h126d:data=8'hFF;
14'h126e:data=8'hFF;
14'h126f:data=8'hFF;
14'h1270:data=8'hFF;
14'h1271:data=8'hFF;
14'h1272:data=8'hC7;
14'h1273:data=8'hC0;
14'h1274:data=8'hC0;
14'h1275:data=8'hC0;
14'h1276:data=8'h00;
14'h1277:data=8'h00;
14'h1278:data=8'h00;
14'h1279:data=8'h00;
14'h127a:data=8'h00;
14'h127b:data=8'h00;
14'h127c:data=8'h00;
14'h127d:data=8'h00;
14'h127e:data=8'h00;
14'h127f:data=8'h00;
14'h1a00:data=8'h00;
14'h1a01:data=8'h00;
14'h1a02:data=8'h00;
14'h1a03:data=8'h00;
14'h1a04:data=8'h00;
14'h1a05:data=8'h00;
14'h1a06:data=8'h00;
14'h1a07:data=8'h00;
14'h1a08:data=8'h00;
14'h1a09:data=8'h00;
14'h1a0a:data=8'h00;
14'h1a0b:data=8'h00;
14'h1a0c:data=8'h00;
14'h1a0d:data=8'h00;
14'h1a0e:data=8'hF8;
14'h1a0f:data=8'hFF;
14'h1a10:data=8'hFF;
14'h1a11:data=8'hFF;
14'h1a12:data=8'hFF;
14'h1a13:data=8'hFF;
14'h1a14:data=8'hFF;
14'h1a15:data=8'hFF;
14'h1a16:data=8'h3F;
14'h1a17:data=8'h01;
14'h1a18:data=8'h00;
14'h1a19:data=8'h00;
14'h1a1a:data=8'h00;
14'h1a1b:data=8'h00;
14'h1a1c:data=8'h00;
14'h1a1d:data=8'h00;
14'h1a1e:data=8'h00;
14'h1a1f:data=8'h00;
14'h1a20:data=8'h00;
14'h1a21:data=8'hC0;
14'h1a22:data=8'hF0;
14'h1a23:data=8'hFC;
14'h1a24:data=8'hFE;
14'h1a25:data=8'hFF;
14'h1a26:data=8'hFF;
14'h1a27:data=8'hFF;
14'h1a28:data=8'hFF;
14'h1a29:data=8'hFF;
14'h1a2a:data=8'h7F;
14'h1a2b:data=8'h3F;
14'h1a2c:data=8'h3F;
14'h1a2d:data=8'h1F;
14'h1a2e:data=8'h3F;
14'h1a2f:data=8'hFF;
14'h1a30:data=8'hFF;
14'h1a31:data=8'hFF;
14'h1a32:data=8'hFF;
14'h1a33:data=8'hFF;
14'h1a34:data=8'hFF;
14'h1a35:data=8'hFF;
14'h1a36:data=8'hFE;
14'h1a37:data=8'hF0;
14'h1a38:data=8'h00;
14'h1a39:data=8'hC0;
14'h1a3a:data=8'hF0;
14'h1a3b:data=8'hF8;
14'h1a3c:data=8'hFE;
14'h1a3d:data=8'hFE;
14'h1a3e:data=8'hFF;
14'h1a3f:data=8'hFF;
14'h1a40:data=8'hFF;
14'h1a41:data=8'hFF;
14'h1a42:data=8'hFF;
14'h1a43:data=8'h7F;
14'h1a44:data=8'h3F;
14'h1a45:data=8'h3F;
14'h1a46:data=8'h1F;
14'h1a47:data=8'h3F;
14'h1a48:data=8'h3F;
14'h1a49:data=8'h3F;
14'h1a4a:data=8'h3F;
14'h1a4b:data=8'h7F;
14'h1a4c:data=8'h07;
14'h1a4d:data=8'hE0;
14'h1a4e:data=8'hF8;
14'h1a4f:data=8'hFC;
14'h1a50:data=8'hFE;
14'h1a51:data=8'hFF;
14'h1a52:data=8'hFF;
14'h1a53:data=8'hFF;
14'h1a54:data=8'hFF;
14'h1a55:data=8'hFF;
14'h1a56:data=8'h7F;
14'h1a57:data=8'h7F;
14'h1a58:data=8'h3F;
14'h1a59:data=8'h3F;
14'h1a5a:data=8'h1F;
14'h1a5b:data=8'hFF;
14'h1a5c:data=8'hFF;
14'h1a5d:data=8'hFF;
14'h1a5e:data=8'hFF;
14'h1a5f:data=8'hFF;
14'h1a60:data=8'hFF;
14'h1a61:data=8'hFF;
14'h1a62:data=8'hFF;
14'h1a63:data=8'h7F;
14'h1a64:data=8'h03;
14'h1a65:data=8'h1F;
14'h1a66:data=8'h1F;
14'h1a67:data=8'hDF;
14'h1a68:data=8'hFF;
14'h1a69:data=8'hFF;
14'h1a6a:data=8'hFF;
14'h1a6b:data=8'hFF;
14'h1a6c:data=8'hFF;
14'h1a6d:data=8'hFF;
14'h1a6e:data=8'hFF;
14'h1a6f:data=8'hFF;
14'h1a70:data=8'h1F;
14'h1a71:data=8'h1F;
14'h1a72:data=8'h1F;
14'h1a73:data=8'h1F;
14'h1a74:data=8'h1F;
14'h1a75:data=8'h0F;
14'h1a76:data=8'h00;
14'h1a77:data=8'h00;
14'h1a78:data=8'h00;
14'h1a79:data=8'h00;
14'h1a7a:data=8'h00;
14'h1a7b:data=8'h00;
14'h1a7c:data=8'h00;
14'h1a7d:data=8'h00;
14'h1a7e:data=8'h00;
14'h1a7f:data=8'h00;
14'h2200:data=8'h00;
14'h2201:data=8'h00;
14'h2202:data=8'h00;
14'h2203:data=8'h00;
14'h2204:data=8'h00;
14'h2205:data=8'h00;
14'h2206:data=8'h00;
14'h2207:data=8'h00;
14'h2208:data=8'h00;
14'h2209:data=8'h00;
14'h220a:data=8'h00;
14'h220b:data=8'h00;
14'h220c:data=8'hF0;
14'h220d:data=8'hFF;
14'h220e:data=8'hFF;
14'h220f:data=8'hFF;
14'h2210:data=8'hFF;
14'h2211:data=8'hFF;
14'h2212:data=8'hFF;
14'h2213:data=8'hFF;
14'h2214:data=8'hFF;
14'h2215:data=8'h87;
14'h2216:data=8'h80;
14'h2217:data=8'h80;
14'h2218:data=8'h80;
14'h2219:data=8'h80;
14'h221a:data=8'h80;
14'h221b:data=8'h80;
14'h221c:data=8'h80;
14'h221d:data=8'h80;
14'h221e:data=8'h80;
14'h221f:data=8'h00;
14'h2220:data=8'h3C;
14'h2221:data=8'hFF;
14'h2222:data=8'hFF;
14'h2223:data=8'hFF;
14'h2224:data=8'hFF;
14'h2225:data=8'hFF;
14'h2226:data=8'hFF;
14'h2227:data=8'hFF;
14'h2228:data=8'hFF;
14'h2229:data=8'hC1;
14'h222a:data=8'hC0;
14'h222b:data=8'h80;
14'h222c:data=8'hC0;
14'h222d:data=8'hE0;
14'h222e:data=8'hF0;
14'h222f:data=8'hFF;
14'h2230:data=8'hFF;
14'h2231:data=8'hFF;
14'h2232:data=8'hFF;
14'h2233:data=8'hFF;
14'h2234:data=8'hFF;
14'h2235:data=8'hFF;
14'h2236:data=8'h7F;
14'h2237:data=8'h0F;
14'h2238:data=8'h00;
14'h2239:data=8'hFF;
14'h223a:data=8'hFF;
14'h223b:data=8'hFF;
14'h223c:data=8'hFF;
14'h223d:data=8'hFF;
14'h223e:data=8'hFF;
14'h223f:data=8'hFF;
14'h2240:data=8'hFF;
14'h2241:data=8'hE3;
14'h2242:data=8'hC0;
14'h2243:data=8'hC0;
14'h2244:data=8'hC0;
14'h2245:data=8'hC0;
14'h2246:data=8'hC0;
14'h2247:data=8'hE0;
14'h2248:data=8'hE0;
14'h2249:data=8'hF0;
14'h224a:data=8'h00;
14'h224b:data=8'h00;
14'h224c:data=8'hFF;
14'h224d:data=8'hFF;
14'h224e:data=8'hFF;
14'h224f:data=8'hFF;
14'h2250:data=8'hFF;
14'h2251:data=8'hFF;
14'h2252:data=8'hFF;
14'h2253:data=8'hFF;
14'h2254:data=8'hE7;
14'h2255:data=8'hC1;
14'h2256:data=8'hC0;
14'h2257:data=8'hC0;
14'h2258:data=8'hE0;
14'h2259:data=8'hF8;
14'h225a:data=8'hFF;
14'h225b:data=8'hFF;
14'h225c:data=8'hFF;
14'h225d:data=8'hFF;
14'h225e:data=8'hFF;
14'h225f:data=8'hFF;
14'h2260:data=8'hFF;
14'h2261:data=8'hFF;
14'h2262:data=8'h0F;
14'h2263:data=8'h00;
14'h2264:data=8'h00;
14'h2265:data=8'h00;
14'h2266:data=8'hF8;
14'h2267:data=8'hFF;
14'h2268:data=8'hFF;
14'h2269:data=8'hFF;
14'h226a:data=8'hFF;
14'h226b:data=8'hFF;
14'h226c:data=8'hFF;
14'h226d:data=8'hFF;
14'h226e:data=8'hFF;
14'h226f:data=8'hC3;
14'h2270:data=8'hC0;
14'h2271:data=8'hE0;
14'h2272:data=8'hE0;
14'h2273:data=8'h00;
14'h2274:data=8'h00;
14'h2275:data=8'h00;
14'h2276:data=8'h00;
14'h2277:data=8'h00;
14'h2278:data=8'h00;
14'h2279:data=8'h00;
14'h227a:data=8'h00;
14'h227b:data=8'h00;
14'h227c:data=8'h00;
14'h227d:data=8'h00;
14'h227e:data=8'h00;
14'h227f:data=8'h00;
14'h2a00:data=8'h00;
14'h2a01:data=8'h00;
14'h2a02:data=8'h00;
14'h2a03:data=8'h00;
14'h2a04:data=8'h00;
14'h2a05:data=8'h00;
14'h2a06:data=8'h00;
14'h2a07:data=8'h00;
14'h2a08:data=8'h00;
14'h2a09:data=8'h00;
14'h2a0a:data=8'h00;
14'h2a0b:data=8'h00;
14'h2a0c:data=8'h1F;
14'h2a0d:data=8'h1F;
14'h2a0e:data=8'h1F;
14'h2a0f:data=8'h1F;
14'h2a10:data=8'h1F;
14'h2a11:data=8'h1F;
14'h2a12:data=8'h1F;
14'h2a13:data=8'h1F;
14'h2a14:data=8'h1F;
14'h2a15:data=8'h1F;
14'h2a16:data=8'h1F;
14'h2a17:data=8'h1F;
14'h2a18:data=8'h1F;
14'h2a19:data=8'h1F;
14'h2a1a:data=8'h1F;
14'h2a1b:data=8'h1F;
14'h2a1c:data=8'h1F;
14'h2a1d:data=8'h1F;
14'h2a1e:data=8'h07;
14'h2a1f:data=8'h00;
14'h2a20:data=8'h00;
14'h2a21:data=8'h01;
14'h2a22:data=8'h07;
14'h2a23:data=8'h0F;
14'h2a24:data=8'h0F;
14'h2a25:data=8'h1F;
14'h2a26:data=8'h1F;
14'h2a27:data=8'h1F;
14'h2a28:data=8'h1F;
14'h2a29:data=8'h1F;
14'h2a2a:data=8'h1F;
14'h2a2b:data=8'h1F;
14'h2a2c:data=8'h1F;
14'h2a2d:data=8'h1F;
14'h2a2e:data=8'h1F;
14'h2a2f:data=8'h1F;
14'h2a30:data=8'h0F;
14'h2a31:data=8'h0F;
14'h2a32:data=8'h07;
14'h2a33:data=8'h07;
14'h2a34:data=8'h03;
14'h2a35:data=8'h01;
14'h2a36:data=8'h00;
14'h2a37:data=8'h00;
14'h2a38:data=8'h00;
14'h2a39:data=8'h01;
14'h2a3a:data=8'h07;
14'h2a3b:data=8'h0F;
14'h2a3c:data=8'h0F;
14'h2a3d:data=8'h1F;
14'h2a3e:data=8'h1F;
14'h2a3f:data=8'h1F;
14'h2a40:data=8'h1F;
14'h2a41:data=8'h1F;
14'h2a42:data=8'h1F;
14'h2a43:data=8'h1F;
14'h2a44:data=8'h1F;
14'h2a45:data=8'h1F;
14'h2a46:data=8'h1F;
14'h2a47:data=8'h0F;
14'h2a48:data=8'h0F;
14'h2a49:data=8'h01;
14'h2a4a:data=8'h00;
14'h2a4b:data=8'h00;
14'h2a4c:data=8'h01;
14'h2a4d:data=8'h07;
14'h2a4e:data=8'h0F;
14'h2a4f:data=8'h1F;
14'h2a50:data=8'h1F;
14'h2a51:data=8'h1F;
14'h2a52:data=8'h1F;
14'h2a53:data=8'h1F;
14'h2a54:data=8'h1F;
14'h2a55:data=8'h1F;
14'h2a56:data=8'h1F;
14'h2a57:data=8'h0F;
14'h2a58:data=8'h0F;
14'h2a59:data=8'h1F;
14'h2a5a:data=8'h1F;
14'h2a5b:data=8'h1F;
14'h2a5c:data=8'h1F;
14'h2a5d:data=8'h1F;
14'h2a5e:data=8'h1F;
14'h2a5f:data=8'h1F;
14'h2a60:data=8'h1F;
14'h2a61:data=8'h01;
14'h2a62:data=8'h00;
14'h2a63:data=8'h00;
14'h2a64:data=8'h00;
14'h2a65:data=8'h00;
14'h2a66:data=8'h07;
14'h2a67:data=8'h0F;
14'h2a68:data=8'h1F;
14'h2a69:data=8'h1F;
14'h2a6a:data=8'h1F;
14'h2a6b:data=8'h1F;
14'h2a6c:data=8'h1F;
14'h2a6d:data=8'h1F;
14'h2a6e:data=8'h1F;
14'h2a6f:data=8'h1F;
14'h2a70:data=8'h1F;
14'h2a71:data=8'h1F;
14'h2a72:data=8'h01;
14'h2a73:data=8'h00;
14'h2a74:data=8'h00;
14'h2a75:data=8'h00;
14'h2a76:data=8'h00;
14'h2a77:data=8'h00;
14'h2a78:data=8'h00;
14'h2a79:data=8'h00;
14'h2a7a:data=8'h00;
14'h2a7b:data=8'h00;
14'h2a7c:data=8'h00;
14'h2a7d:data=8'h00;
14'h2a7e:data=8'h00;
14'h2a7f:data=8'h00;
14'h3200:data=8'h00;
14'h3201:data=8'h00;
14'h3202:data=8'h00;
14'h3203:data=8'h00;
14'h3204:data=8'h00;
14'h3205:data=8'h00;
14'h3206:data=8'h00;
14'h3207:data=8'h00;
14'h3208:data=8'h00;
14'h3209:data=8'h00;
14'h320a:data=8'h00;
14'h320b:data=8'h00;
14'h320c:data=8'h00;
14'h320d:data=8'h00;
14'h320e:data=8'h00;
14'h320f:data=8'h00;
14'h3210:data=8'h00;
14'h3211:data=8'h00;
14'h3212:data=8'h00;
14'h3213:data=8'h00;
14'h3214:data=8'h00;
14'h3215:data=8'h00;
14'h3216:data=8'h00;
14'h3217:data=8'h00;
14'h3218:data=8'h00;
14'h3219:data=8'h00;
14'h321a:data=8'h00;
14'h321b:data=8'h00;
14'h321c:data=8'h00;
14'h321d:data=8'h00;
14'h321e:data=8'h00;
14'h321f:data=8'h00;
14'h3220:data=8'h00;
14'h3221:data=8'h00;
14'h3222:data=8'h00;
14'h3223:data=8'h00;
14'h3224:data=8'h00;
14'h3225:data=8'h00;
14'h3226:data=8'h00;
14'h3227:data=8'h00;
14'h3228:data=8'h00;
14'h3229:data=8'h00;
14'h322a:data=8'h00;
14'h322b:data=8'h00;
14'h322c:data=8'h00;
14'h322d:data=8'h00;
14'h322e:data=8'h00;
14'h322f:data=8'h00;
14'h3230:data=8'h00;
14'h3231:data=8'h00;
14'h3232:data=8'h00;
14'h3233:data=8'h00;
14'h3234:data=8'h00;
14'h3235:data=8'h00;
14'h3236:data=8'h00;
14'h3237:data=8'h00;
14'h3238:data=8'h00;
14'h3239:data=8'h00;
14'h323a:data=8'h00;
14'h323b:data=8'h00;
14'h323c:data=8'h00;
14'h323d:data=8'h00;
14'h323e:data=8'h00;
14'h323f:data=8'h00;
14'h3240:data=8'h00;
14'h3241:data=8'h00;
14'h3242:data=8'h00;
14'h3243:data=8'h00;
14'h3244:data=8'h00;
14'h3245:data=8'h00;
14'h3246:data=8'h00;
14'h3247:data=8'h00;
14'h3248:data=8'h00;
14'h3249:data=8'h00;
14'h324a:data=8'h00;
14'h324b:data=8'h00;
14'h324c:data=8'h00;
14'h324d:data=8'h00;
14'h324e:data=8'h00;
14'h324f:data=8'h00;
14'h3250:data=8'h00;
14'h3251:data=8'h00;
14'h3252:data=8'h00;
14'h3253:data=8'h00;
14'h3254:data=8'h00;
14'h3255:data=8'h00;
14'h3256:data=8'h00;
14'h3257:data=8'h00;
14'h3258:data=8'h00;
14'h3259:data=8'h00;
14'h325a:data=8'h00;
14'h325b:data=8'h00;
14'h325c:data=8'h00;
14'h325d:data=8'h00;
14'h325e:data=8'h00;
14'h325f:data=8'h00;
14'h3260:data=8'h00;
14'h3261:data=8'h00;
14'h3262:data=8'h00;
14'h3263:data=8'h00;
14'h3264:data=8'h00;
14'h3265:data=8'h00;
14'h3266:data=8'h00;
14'h3267:data=8'h00;
14'h3268:data=8'h00;
14'h3269:data=8'h00;
14'h326a:data=8'h00;
14'h326b:data=8'h00;
14'h326c:data=8'h00;
14'h326d:data=8'h00;
14'h326e:data=8'h00;
14'h326f:data=8'h00;
14'h3270:data=8'h00;
14'h3271:data=8'h00;
14'h3272:data=8'h00;
14'h3273:data=8'h00;
14'h3274:data=8'h00;
14'h3275:data=8'h00;
14'h3276:data=8'h00;
14'h3277:data=8'h00;
14'h3278:data=8'h00;
14'h3279:data=8'h00;
14'h327a:data=8'h00;
14'h327b:data=8'h00;
14'h327c:data=8'h00;
14'h327d:data=8'h00;
14'h327e:data=8'h00;
14'h327f:data=8'h00;
14'h3a00:data=8'h00;
14'h3a01:data=8'h00;
14'h3a02:data=8'h00;
14'h3a03:data=8'h00;
14'h3a04:data=8'h00;
14'h3a05:data=8'h00;
14'h3a06:data=8'h00;
14'h3a07:data=8'h00;
14'h3a08:data=8'h00;
14'h3a09:data=8'h00;
14'h3a0a:data=8'h00;
14'h3a0b:data=8'h00;
14'h3a0c:data=8'h00;
14'h3a0d:data=8'h00;
14'h3a0e:data=8'h00;
14'h3a0f:data=8'h00;
14'h3a10:data=8'h00;
14'h3a11:data=8'h00;
14'h3a12:data=8'h00;
14'h3a13:data=8'h00;
14'h3a14:data=8'h00;
14'h3a15:data=8'h00;
14'h3a16:data=8'h00;
14'h3a17:data=8'h00;
14'h3a18:data=8'h00;
14'h3a19:data=8'h00;
14'h3a1a:data=8'h00;
14'h3a1b:data=8'h00;
14'h3a1c:data=8'h00;
14'h3a1d:data=8'h00;
14'h3a1e:data=8'h00;
14'h3a1f:data=8'h00;
14'h3a20:data=8'h00;
14'h3a21:data=8'h00;
14'h3a22:data=8'h00;
14'h3a23:data=8'h00;
14'h3a24:data=8'h00;
14'h3a25:data=8'h00;
14'h3a26:data=8'h00;
14'h3a27:data=8'h00;
14'h3a28:data=8'h00;
14'h3a29:data=8'h00;
14'h3a2a:data=8'h00;
14'h3a2b:data=8'h00;
14'h3a2c:data=8'h00;
14'h3a2d:data=8'h00;
14'h3a2e:data=8'h00;
14'h3a2f:data=8'h00;
14'h3a30:data=8'h00;
14'h3a31:data=8'h00;
14'h3a32:data=8'h00;
14'h3a33:data=8'h00;
14'h3a34:data=8'h00;
14'h3a35:data=8'h00;
14'h3a36:data=8'h00;
14'h3a37:data=8'h00;
14'h3a38:data=8'h00;
14'h3a39:data=8'h00;
14'h3a3a:data=8'h00;
14'h3a3b:data=8'h00;
14'h3a3c:data=8'h00;
14'h3a3d:data=8'h00;
14'h3a3e:data=8'h00;
14'h3a3f:data=8'h00;
14'h3a40:data=8'h00;
14'h3a41:data=8'h00;
14'h3a42:data=8'h00;
14'h3a43:data=8'h00;
14'h3a44:data=8'h00;
14'h3a45:data=8'h00;
14'h3a46:data=8'h00;
14'h3a47:data=8'h00;
14'h3a48:data=8'h00;
14'h3a49:data=8'h00;
14'h3a4a:data=8'h00;
14'h3a4b:data=8'h00;
14'h3a4c:data=8'h00;
14'h3a4d:data=8'h00;
14'h3a4e:data=8'h00;
14'h3a4f:data=8'h00;
14'h3a50:data=8'h00;
14'h3a51:data=8'h00;
14'h3a52:data=8'h00;
14'h3a53:data=8'h00;
14'h3a54:data=8'h00;
14'h3a55:data=8'h00;
14'h3a56:data=8'h00;
14'h3a57:data=8'h00;
14'h3a58:data=8'h00;
14'h3a59:data=8'h00;
14'h3a5a:data=8'h00;
14'h3a5b:data=8'h00;
14'h3a5c:data=8'h00;
14'h3a5d:data=8'h00;
14'h3a5e:data=8'h00;
14'h3a5f:data=8'h00;
14'h3a60:data=8'h00;
14'h3a61:data=8'h00;
14'h3a62:data=8'h00;
14'h3a63:data=8'h00;
14'h3a64:data=8'h00;
14'h3a65:data=8'h00;
14'h3a66:data=8'h00;
14'h3a67:data=8'h00;
14'h3a68:data=8'h00;
14'h3a69:data=8'h00;
14'h3a6a:data=8'h00;
14'h3a6b:data=8'h00;
14'h3a6c:data=8'h00;
14'h3a6d:data=8'h00;
14'h3a6e:data=8'h00;
14'h3a6f:data=8'h00;
14'h3a70:data=8'h00;
14'h3a71:data=8'h00;
14'h3a72:data=8'h00;
14'h3a73:data=8'h00;
14'h3a74:data=8'h00;
14'h3a75:data=8'h00;
14'h3a76:data=8'h00;
14'h3a77:data=8'h00;
14'h3a78:data=8'h00;
14'h3a79:data=8'h00;
14'h3a7a:data=8'h00;
14'h3a7b:data=8'h00;
14'h3a7c:data=8'h00;
14'h3a7d:data=8'h00;
14'h3a7e:data=8'h00;
14'h3a7f:data=8'h00;
///////////////////////////////////////////////////////////////////////////PIC4 Light
14'h0300:data=8'h00;
14'h0301:data=8'h00;
14'h0302:data=8'h00;
14'h0303:data=8'h00;
14'h0304:data=8'h00;
14'h0305:data=8'h00;
14'h0306:data=8'h00;
14'h0307:data=8'h00;
14'h0308:data=8'h00;
14'h0309:data=8'h00;
14'h030a:data=8'h00;
14'h030b:data=8'h00;
14'h030c:data=8'h00;
14'h030d:data=8'h00;
14'h030e:data=8'h00;
14'h030f:data=8'h00;
14'h0310:data=8'h00;
14'h0311:data=8'h00;
14'h0312:data=8'h00;
14'h0313:data=8'h00;
14'h0314:data=8'h00;
14'h0315:data=8'h00;
14'h0316:data=8'h00;
14'h0317:data=8'h00;
14'h0318:data=8'h00;
14'h0319:data=8'h00;
14'h031a:data=8'h00;
14'h031b:data=8'h00;
14'h031c:data=8'h00;
14'h031d:data=8'h00;
14'h031e:data=8'h00;
14'h031f:data=8'h00;
14'h0320:data=8'h00;
14'h0321:data=8'h00;
14'h0322:data=8'h00;
14'h0323:data=8'h00;
14'h0324:data=8'h00;
14'h0325:data=8'h00;
14'h0326:data=8'h00;
14'h0327:data=8'h00;
14'h0328:data=8'h00;
14'h0329:data=8'h00;
14'h032a:data=8'h00;
14'h032b:data=8'h00;
14'h032c:data=8'h00;
14'h032d:data=8'h00;
14'h032e:data=8'h00;
14'h032f:data=8'h00;
14'h0330:data=8'h00;
14'h0331:data=8'h00;
14'h0332:data=8'h00;
14'h0333:data=8'h00;
14'h0334:data=8'h00;
14'h0335:data=8'h00;
14'h0336:data=8'h00;
14'h0337:data=8'h00;
14'h0338:data=8'h00;
14'h0339:data=8'h00;
14'h033a:data=8'h00;
14'h033b:data=8'h00;
14'h033c:data=8'h00;
14'h033d:data=8'h00;
14'h033e:data=8'h00;
14'h033f:data=8'h00;
14'h0340:data=8'h00;
14'h0341:data=8'h00;
14'h0342:data=8'h00;
14'h0343:data=8'h00;
14'h0344:data=8'h00;
14'h0345:data=8'h00;
14'h0346:data=8'h00;
14'h0347:data=8'h00;
14'h0348:data=8'h00;
14'h0349:data=8'h00;
14'h034a:data=8'h00;
14'h034b:data=8'h00;
14'h034c:data=8'h00;
14'h034d:data=8'h00;
14'h034e:data=8'h00;
14'h034f:data=8'h00;
14'h0350:data=8'h00;
14'h0351:data=8'h00;
14'h0352:data=8'h00;
14'h0353:data=8'h00;
14'h0354:data=8'h00;
14'h0355:data=8'h00;
14'h0356:data=8'h00;
14'h0357:data=8'h00;
14'h0358:data=8'h00;
14'h0359:data=8'h00;
14'h035a:data=8'h00;
14'h035b:data=8'h00;
14'h035c:data=8'h00;
14'h035d:data=8'h00;
14'h035e:data=8'h00;
14'h035f:data=8'h00;
14'h0360:data=8'h00;
14'h0361:data=8'h00;
14'h0362:data=8'h00;
14'h0363:data=8'h00;
14'h0364:data=8'h00;
14'h0365:data=8'h00;
14'h0366:data=8'h00;
14'h0367:data=8'h00;
14'h0368:data=8'h00;
14'h0369:data=8'h00;
14'h036a:data=8'h00;
14'h036b:data=8'h00;
14'h036c:data=8'h00;
14'h036d:data=8'h00;
14'h036e:data=8'h00;
14'h036f:data=8'h00;
14'h0370:data=8'h00;
14'h0371:data=8'h00;
14'h0372:data=8'h00;
14'h0373:data=8'h00;
14'h0374:data=8'h00;
14'h0375:data=8'h00;
14'h0376:data=8'h00;
14'h0377:data=8'h00;
14'h0378:data=8'h00;
14'h0379:data=8'h00;
14'h037a:data=8'h00;
14'h037b:data=8'h00;
14'h037c:data=8'h00;
14'h037d:data=8'h00;
14'h037e:data=8'h00;
14'h037f:data=8'h00;
14'h0b00:data=8'h00;
14'h0b01:data=8'h00;
14'h0b02:data=8'h00;
14'h0b03:data=8'h00;
14'h0b04:data=8'h00;
14'h0b05:data=8'h00;
14'h0b06:data=8'h00;
14'h0b07:data=8'h00;
14'h0b08:data=8'h00;
14'h0b09:data=8'h00;
14'h0b0a:data=8'h00;
14'h0b0b:data=8'h00;
14'h0b0c:data=8'h00;
14'h0b0d:data=8'h00;
14'h0b0e:data=8'h00;
14'h0b0f:data=8'h00;
14'h0b10:data=8'h00;
14'h0b11:data=8'h00;
14'h0b12:data=8'h00;
14'h0b13:data=8'h00;
14'h0b14:data=8'h00;
14'h0b15:data=8'h00;
14'h0b16:data=8'h00;
14'h0b17:data=8'h00;
14'h0b18:data=8'h00;
14'h0b19:data=8'h00;
14'h0b1a:data=8'h00;
14'h0b1b:data=8'h00;
14'h0b1c:data=8'h00;
14'h0b1d:data=8'h00;
14'h0b1e:data=8'h00;
14'h0b1f:data=8'h00;
14'h0b20:data=8'h00;
14'h0b21:data=8'h00;
14'h0b22:data=8'h00;
14'h0b23:data=8'h00;
14'h0b24:data=8'h00;
14'h0b25:data=8'h00;
14'h0b26:data=8'h00;
14'h0b27:data=8'h80;
14'h0b28:data=8'hC0;
14'h0b29:data=8'hC0;
14'h0b2a:data=8'hC0;
14'h0b2b:data=8'hC0;
14'h0b2c:data=8'hC0;
14'h0b2d:data=8'hC0;
14'h0b2e:data=8'hC0;
14'h0b2f:data=8'h80;
14'h0b30:data=8'h00;
14'h0b31:data=8'h00;
14'h0b32:data=8'h00;
14'h0b33:data=8'h00;
14'h0b34:data=8'h00;
14'h0b35:data=8'h00;
14'h0b36:data=8'h00;
14'h0b37:data=8'h00;
14'h0b38:data=8'h00;
14'h0b39:data=8'h00;
14'h0b3a:data=8'h00;
14'h0b3b:data=8'h00;
14'h0b3c:data=8'h00;
14'h0b3d:data=8'h00;
14'h0b3e:data=8'h00;
14'h0b3f:data=8'h00;
14'h0b40:data=8'h00;
14'h0b41:data=8'h00;
14'h0b42:data=8'h00;
14'h0b43:data=8'h00;
14'h0b44:data=8'h00;
14'h0b45:data=8'h00;
14'h0b46:data=8'h00;
14'h0b47:data=8'h00;
14'h0b48:data=8'h00;
14'h0b49:data=8'h00;
14'h0b4a:data=8'h00;
14'h0b4b:data=8'h00;
14'h0b4c:data=8'h00;
14'h0b4d:data=8'h00;
14'h0b4e:data=8'hC0;
14'h0b4f:data=8'hC0;
14'h0b50:data=8'hC0;
14'h0b51:data=8'hC0;
14'h0b52:data=8'hC0;
14'h0b53:data=8'hC0;
14'h0b54:data=8'hC0;
14'h0b55:data=8'hC0;
14'h0b56:data=8'hC0;
14'h0b57:data=8'h00;
14'h0b58:data=8'h00;
14'h0b59:data=8'h00;
14'h0b5a:data=8'h00;
14'h0b5b:data=8'h00;
14'h0b5c:data=8'h00;
14'h0b5d:data=8'h00;
14'h0b5e:data=8'h00;
14'h0b5f:data=8'h00;
14'h0b60:data=8'h00;
14'h0b61:data=8'h00;
14'h0b62:data=8'h00;
14'h0b63:data=8'h00;
14'h0b64:data=8'h00;
14'h0b65:data=8'h00;
14'h0b66:data=8'h00;
14'h0b67:data=8'h00;
14'h0b68:data=8'h00;
14'h0b69:data=8'h00;
14'h0b6a:data=8'h00;
14'h0b6b:data=8'h00;
14'h0b6c:data=8'h00;
14'h0b6d:data=8'h00;
14'h0b6e:data=8'h00;
14'h0b6f:data=8'h00;
14'h0b70:data=8'h00;
14'h0b71:data=8'h00;
14'h0b72:data=8'h00;
14'h0b73:data=8'h00;
14'h0b74:data=8'h00;
14'h0b75:data=8'h00;
14'h0b76:data=8'h00;
14'h0b77:data=8'h00;
14'h0b78:data=8'h00;
14'h0b79:data=8'h00;
14'h0b7a:data=8'h00;
14'h0b7b:data=8'h00;
14'h0b7c:data=8'h00;
14'h0b7d:data=8'h00;
14'h0b7e:data=8'h00;
14'h0b7f:data=8'h00;
14'h1300:data=8'h00;
14'h1301:data=8'h00;
14'h1302:data=8'h00;
14'h1303:data=8'h00;
14'h1304:data=8'h00;
14'h1305:data=8'h00;
14'h1306:data=8'h00;
14'h1307:data=8'h00;
14'h1308:data=8'h00;
14'h1309:data=8'h00;
14'h130a:data=8'h00;
14'h130b:data=8'h00;
14'h130c:data=8'h00;
14'h130d:data=8'h00;
14'h130e:data=8'h00;
14'h130f:data=8'h00;
14'h1310:data=8'h00;
14'h1311:data=8'hC0;
14'h1312:data=8'hFC;
14'h1313:data=8'hFF;
14'h1314:data=8'hFF;
14'h1315:data=8'hFF;
14'h1316:data=8'hFF;
14'h1317:data=8'hFF;
14'h1318:data=8'hFF;
14'h1319:data=8'hFF;
14'h131a:data=8'h3F;
14'h131b:data=8'h00;
14'h131c:data=8'h00;
14'h131d:data=8'h00;
14'h131e:data=8'h00;
14'h131f:data=8'h00;
14'h1320:data=8'h00;
14'h1321:data=8'h00;
14'h1322:data=8'h00;
14'h1323:data=8'h00;
14'h1324:data=8'h00;
14'h1325:data=8'h00;
14'h1326:data=8'h00;
14'h1327:data=8'h1F;
14'h1328:data=8'h3F;
14'h1329:data=8'h7F;
14'h132a:data=8'h7F;
14'h132b:data=8'h7F;
14'h132c:data=8'h7F;
14'h132d:data=8'h7F;
14'h132e:data=8'h3F;
14'h132f:data=8'h1F;
14'h1330:data=8'h00;
14'h1331:data=8'h00;
14'h1332:data=8'h00;
14'h1333:data=8'h00;
14'h1334:data=8'h00;
14'h1335:data=8'h00;
14'h1336:data=8'h00;
14'h1337:data=8'h00;
14'h1338:data=8'h00;
14'h1339:data=8'h00;
14'h133a:data=8'h00;
14'h133b:data=8'h00;
14'h133c:data=8'h00;
14'h133d:data=8'h00;
14'h133e:data=8'h00;
14'h133f:data=8'h00;
14'h1340:data=8'h00;
14'h1341:data=8'h00;
14'h1342:data=8'h00;
14'h1343:data=8'h00;
14'h1344:data=8'h00;
14'h1345:data=8'h00;
14'h1346:data=8'h00;
14'h1347:data=8'h00;
14'h1348:data=8'h00;
14'h1349:data=8'h00;
14'h134a:data=8'h00;
14'h134b:data=8'h00;
14'h134c:data=8'hC0;
14'h134d:data=8'hFC;
14'h134e:data=8'hFF;
14'h134f:data=8'hFF;
14'h1350:data=8'hFF;
14'h1351:data=8'hFF;
14'h1352:data=8'hFF;
14'h1353:data=8'hFF;
14'h1354:data=8'hFF;
14'h1355:data=8'h1F;
14'h1356:data=8'h01;
14'h1357:data=8'h00;
14'h1358:data=8'h00;
14'h1359:data=8'h00;
14'h135a:data=8'h00;
14'h135b:data=8'h00;
14'h135c:data=8'h00;
14'h135d:data=8'h00;
14'h135e:data=8'h00;
14'h135f:data=8'h00;
14'h1360:data=8'h00;
14'h1361:data=8'h00;
14'h1362:data=8'h00;
14'h1363:data=8'h00;
14'h1364:data=8'h00;
14'h1365:data=8'h00;
14'h1366:data=8'hE0;
14'h1367:data=8'hFC;
14'h1368:data=8'hFC;
14'h1369:data=8'hFC;
14'h136a:data=8'hFE;
14'h136b:data=8'hFE;
14'h136c:data=8'hFE;
14'h136d:data=8'hFE;
14'h136e:data=8'hFE;
14'h136f:data=8'h06;
14'h1370:data=8'h00;
14'h1371:data=8'h00;
14'h1372:data=8'h00;
14'h1373:data=8'h00;
14'h1374:data=8'h00;
14'h1375:data=8'h00;
14'h1376:data=8'h00;
14'h1377:data=8'h00;
14'h1378:data=8'h00;
14'h1379:data=8'h00;
14'h137a:data=8'h00;
14'h137b:data=8'h00;
14'h137c:data=8'h00;
14'h137d:data=8'h00;
14'h137e:data=8'h00;
14'h137f:data=8'h00;
14'h1b00:data=8'h00;
14'h1b01:data=8'h00;
14'h1b02:data=8'h00;
14'h1b03:data=8'h00;
14'h1b04:data=8'h00;
14'h1b05:data=8'h00;
14'h1b06:data=8'h00;
14'h1b07:data=8'h00;
14'h1b08:data=8'h00;
14'h1b09:data=8'h00;
14'h1b0a:data=8'h00;
14'h1b0b:data=8'h00;
14'h1b0c:data=8'h00;
14'h1b0d:data=8'h00;
14'h1b0e:data=8'h00;
14'h1b0f:data=8'h00;
14'h1b10:data=8'hF8;
14'h1b11:data=8'hFF;
14'h1b12:data=8'hFF;
14'h1b13:data=8'hFF;
14'h1b14:data=8'hFF;
14'h1b15:data=8'hFF;
14'h1b16:data=8'hFF;
14'h1b17:data=8'hFF;
14'h1b18:data=8'hFF;
14'h1b19:data=8'h07;
14'h1b1a:data=8'h00;
14'h1b1b:data=8'h00;
14'h1b1c:data=8'h00;
14'h1b1d:data=8'h00;
14'h1b1e:data=8'h00;
14'h1b1f:data=8'h00;
14'h1b20:data=8'h00;
14'h1b21:data=8'h00;
14'h1b22:data=8'h00;
14'h1b23:data=8'h00;
14'h1b24:data=8'hC0;
14'h1b25:data=8'hFC;
14'h1b26:data=8'hFF;
14'h1b27:data=8'hFF;
14'h1b28:data=8'hFF;
14'h1b29:data=8'hFF;
14'h1b2a:data=8'hFF;
14'h1b2b:data=8'hFF;
14'h1b2c:data=8'hFF;
14'h1b2d:data=8'h1F;
14'h1b2e:data=8'h00;
14'h1b2f:data=8'h00;
14'h1b30:data=8'h00;
14'h1b31:data=8'hC0;
14'h1b32:data=8'hE0;
14'h1b33:data=8'hF0;
14'h1b34:data=8'hF8;
14'h1b35:data=8'hFC;
14'h1b36:data=8'hFE;
14'h1b37:data=8'hFE;
14'h1b38:data=8'hFF;
14'h1b39:data=8'hFF;
14'h1b3a:data=8'hFF;
14'h1b3b:data=8'hFF;
14'h1b3c:data=8'hFF;
14'h1b3d:data=8'h7F;
14'h1b3e:data=8'h7F;
14'h1b3f:data=8'hFF;
14'h1b40:data=8'hFF;
14'h1b41:data=8'hFF;
14'h1b42:data=8'hFF;
14'h1b43:data=8'hFF;
14'h1b44:data=8'hFF;
14'h1b45:data=8'hFF;
14'h1b46:data=8'hFF;
14'h1b47:data=8'h7E;
14'h1b48:data=8'h00;
14'h1b49:data=8'h00;
14'h1b4a:data=8'h00;
14'h1b4b:data=8'hF8;
14'h1b4c:data=8'hFF;
14'h1b4d:data=8'hFF;
14'h1b4e:data=8'hFF;
14'h1b4f:data=8'hFF;
14'h1b50:data=8'hFF;
14'h1b51:data=8'hFF;
14'h1b52:data=8'hFF;
14'h1b53:data=8'hFF;
14'h1b54:data=8'hFF;
14'h1b55:data=8'hFE;
14'h1b56:data=8'hFF;
14'h1b57:data=8'h7F;
14'h1b58:data=8'hFF;
14'h1b59:data=8'hFF;
14'h1b5a:data=8'hFF;
14'h1b5b:data=8'hFF;
14'h1b5c:data=8'hFF;
14'h1b5d:data=8'hFF;
14'h1b5e:data=8'hFF;
14'h1b5f:data=8'hFE;
14'h1b60:data=8'hF8;
14'h1b61:data=8'h00;
14'h1b62:data=8'h7E;
14'h1b63:data=8'h7F;
14'h1b64:data=8'hFF;
14'h1b65:data=8'hFF;
14'h1b66:data=8'hFF;
14'h1b67:data=8'hFF;
14'h1b68:data=8'hFF;
14'h1b69:data=8'hFF;
14'h1b6a:data=8'hFF;
14'h1b6b:data=8'hFF;
14'h1b6c:data=8'hFF;
14'h1b6d:data=8'h7F;
14'h1b6e:data=8'h7F;
14'h1b6f:data=8'h7F;
14'h1b70:data=8'h7F;
14'h1b71:data=8'h7F;
14'h1b72:data=8'h1F;
14'h1b73:data=8'h00;
14'h1b74:data=8'h00;
14'h1b75:data=8'h00;
14'h1b76:data=8'h00;
14'h1b77:data=8'h00;
14'h1b78:data=8'h00;
14'h1b79:data=8'h00;
14'h1b7a:data=8'h00;
14'h1b7b:data=8'h00;
14'h1b7c:data=8'h00;
14'h1b7d:data=8'h00;
14'h1b7e:data=8'h00;
14'h1b7f:data=8'h00;
14'h2300:data=8'h00;
14'h2301:data=8'h00;
14'h2302:data=8'h00;
14'h2303:data=8'h00;
14'h2304:data=8'h00;
14'h2305:data=8'h00;
14'h2306:data=8'h00;
14'h2307:data=8'h00;
14'h2308:data=8'h00;
14'h2309:data=8'h00;
14'h230a:data=8'h00;
14'h230b:data=8'h00;
14'h230c:data=8'h00;
14'h230d:data=8'h00;
14'h230e:data=8'hE0;
14'h230f:data=8'hFF;
14'h2310:data=8'hFF;
14'h2311:data=8'hFF;
14'h2312:data=8'hFF;
14'h2313:data=8'hFF;
14'h2314:data=8'hFF;
14'h2315:data=8'hFF;
14'h2316:data=8'hFF;
14'h2317:data=8'h0F;
14'h2318:data=8'h00;
14'h2319:data=8'h00;
14'h231a:data=8'h00;
14'h231b:data=8'h00;
14'h231c:data=8'h00;
14'h231d:data=8'h00;
14'h231e:data=8'h00;
14'h231f:data=8'h00;
14'h2320:data=8'h00;
14'h2321:data=8'h00;
14'h2322:data=8'h00;
14'h2323:data=8'hF8;
14'h2324:data=8'hFF;
14'h2325:data=8'hFF;
14'h2326:data=8'hFF;
14'h2327:data=8'hFF;
14'h2328:data=8'hFF;
14'h2329:data=8'hFF;
14'h232a:data=8'hFF;
14'h232b:data=8'h7F;
14'h232c:data=8'h03;
14'h232d:data=8'h00;
14'h232e:data=8'h00;
14'h232f:data=8'h00;
14'h2330:data=8'hFF;
14'h2331:data=8'hFF;
14'h2332:data=8'hFF;
14'h2333:data=8'hFF;
14'h2334:data=8'hFF;
14'h2335:data=8'hFF;
14'h2336:data=8'hFF;
14'h2337:data=8'hFF;
14'h2338:data=8'h0F;
14'h2339:data=8'h03;
14'h233a:data=8'h01;
14'h233b:data=8'h80;
14'h233c:data=8'hC0;
14'h233d:data=8'hF0;
14'h233e:data=8'hFE;
14'h233f:data=8'hFF;
14'h2340:data=8'hFF;
14'h2341:data=8'hFF;
14'h2342:data=8'hFF;
14'h2343:data=8'hFF;
14'h2344:data=8'hFF;
14'h2345:data=8'hFF;
14'h2346:data=8'h0F;
14'h2347:data=8'h00;
14'h2348:data=8'h00;
14'h2349:data=8'hE0;
14'h234a:data=8'hFF;
14'h234b:data=8'hFF;
14'h234c:data=8'hFF;
14'h234d:data=8'hFF;
14'h234e:data=8'hFF;
14'h234f:data=8'hFF;
14'h2350:data=8'hFF;
14'h2351:data=8'hFF;
14'h2352:data=8'h0F;
14'h2353:data=8'h03;
14'h2354:data=8'h01;
14'h2355:data=8'h00;
14'h2356:data=8'h00;
14'h2357:data=8'hF8;
14'h2358:data=8'hFF;
14'h2359:data=8'hFF;
14'h235a:data=8'hFF;
14'h235b:data=8'hFF;
14'h235c:data=8'hFF;
14'h235d:data=8'hFF;
14'h235e:data=8'hFF;
14'h235f:data=8'h3F;
14'h2360:data=8'h01;
14'h2361:data=8'h00;
14'h2362:data=8'h00;
14'h2363:data=8'hF8;
14'h2364:data=8'hFF;
14'h2365:data=8'hFF;
14'h2366:data=8'hFF;
14'h2367:data=8'hFF;
14'h2368:data=8'hFF;
14'h2369:data=8'hFF;
14'h236a:data=8'hFF;
14'h236b:data=8'h3F;
14'h236c:data=8'h01;
14'h236d:data=8'h00;
14'h236e:data=8'h80;
14'h236f:data=8'h80;
14'h2370:data=8'h00;
14'h2371:data=8'h00;
14'h2372:data=8'h00;
14'h2373:data=8'h00;
14'h2374:data=8'h00;
14'h2375:data=8'h00;
14'h2376:data=8'h00;
14'h2377:data=8'h00;
14'h2378:data=8'h00;
14'h2379:data=8'h00;
14'h237a:data=8'h00;
14'h237b:data=8'h00;
14'h237c:data=8'h00;
14'h237d:data=8'h00;
14'h237e:data=8'h00;
14'h237f:data=8'h00;
14'h2b00:data=8'h00;
14'h2b01:data=8'h00;
14'h2b02:data=8'h00;
14'h2b03:data=8'h00;
14'h2b04:data=8'h00;
14'h2b05:data=8'h00;
14'h2b06:data=8'h00;
14'h2b07:data=8'h00;
14'h2b08:data=8'h00;
14'h2b09:data=8'h00;
14'h2b0a:data=8'h00;
14'h2b0b:data=8'h00;
14'h2b0c:data=8'h00;
14'h2b0d:data=8'h00;
14'h2b0e:data=8'h7F;
14'h2b0f:data=8'h7F;
14'h2b10:data=8'h7F;
14'h2b11:data=8'h7F;
14'h2b12:data=8'h7F;
14'h2b13:data=8'h7F;
14'h2b14:data=8'h7F;
14'h2b15:data=8'h7F;
14'h2b16:data=8'h7F;
14'h2b17:data=8'h7E;
14'h2b18:data=8'h7E;
14'h2b19:data=8'h7E;
14'h2b1a:data=8'h7E;
14'h2b1b:data=8'h7E;
14'h2b1c:data=8'h7E;
14'h2b1d:data=8'h7E;
14'h2b1e:data=8'h7E;
14'h2b1f:data=8'h7E;
14'h2b20:data=8'h1E;
14'h2b21:data=8'h00;
14'h2b22:data=8'h00;
14'h2b23:data=8'h1F;
14'h2b24:data=8'h3F;
14'h2b25:data=8'h7F;
14'h2b26:data=8'h7F;
14'h2b27:data=8'h7F;
14'h2b28:data=8'h7F;
14'h2b29:data=8'h7F;
14'h2b2a:data=8'h7F;
14'h2b2b:data=8'h7F;
14'h2b2c:data=8'h7F;
14'h2b2d:data=8'h7F;
14'h2b2e:data=8'h0F;
14'h2b2f:data=8'h00;
14'h2b30:data=8'h87;
14'h2b31:data=8'h1F;
14'h2b32:data=8'h3F;
14'h2b33:data=8'h7F;
14'h2b34:data=8'h7F;
14'h2b35:data=8'h7F;
14'h2b36:data=8'h7F;
14'h2b37:data=8'h7F;
14'h2b38:data=8'h7F;
14'h2b39:data=8'h7F;
14'h2b3a:data=8'hFF;
14'h2b3b:data=8'hFF;
14'h2b3c:data=8'hFF;
14'h2b3d:data=8'hFF;
14'h2b3e:data=8'hFF;
14'h2b3f:data=8'hFF;
14'h2b40:data=8'hFF;
14'h2b41:data=8'hFF;
14'h2b42:data=8'hFF;
14'h2b43:data=8'hFF;
14'h2b44:data=8'h1F;
14'h2b45:data=8'h00;
14'h2b46:data=8'h00;
14'h2b47:data=8'h00;
14'h2b48:data=8'h7C;
14'h2b49:data=8'h7F;
14'h2b4a:data=8'h7F;
14'h2b4b:data=8'h7F;
14'h2b4c:data=8'h7F;
14'h2b4d:data=8'h7F;
14'h2b4e:data=8'h7F;
14'h2b4f:data=8'h7F;
14'h2b50:data=8'h1F;
14'h2b51:data=8'h00;
14'h2b52:data=8'h00;
14'h2b53:data=8'h00;
14'h2b54:data=8'h00;
14'h2b55:data=8'h60;
14'h2b56:data=8'h7F;
14'h2b57:data=8'h7F;
14'h2b58:data=8'h7F;
14'h2b59:data=8'h7F;
14'h2b5a:data=8'h7F;
14'h2b5b:data=8'h7F;
14'h2b5c:data=8'h7F;
14'h2b5d:data=8'h7F;
14'h2b5e:data=8'h07;
14'h2b5f:data=8'h00;
14'h2b60:data=8'h00;
14'h2b61:data=8'h00;
14'h2b62:data=8'h00;
14'h2b63:data=8'h1F;
14'h2b64:data=8'h3F;
14'h2b65:data=8'h7F;
14'h2b66:data=8'h7F;
14'h2b67:data=8'h7F;
14'h2b68:data=8'h7F;
14'h2b69:data=8'h7F;
14'h2b6a:data=8'h7F;
14'h2b6b:data=8'h7F;
14'h2b6c:data=8'h7F;
14'h2b6d:data=8'h7F;
14'h2b6e:data=8'h3F;
14'h2b6f:data=8'h03;
14'h2b70:data=8'h00;
14'h2b71:data=8'h00;
14'h2b72:data=8'h00;
14'h2b73:data=8'h00;
14'h2b74:data=8'h00;
14'h2b75:data=8'h00;
14'h2b76:data=8'h00;
14'h2b77:data=8'h00;
14'h2b78:data=8'h00;
14'h2b79:data=8'h00;
14'h2b7a:data=8'h00;
14'h2b7b:data=8'h00;
14'h2b7c:data=8'h00;
14'h2b7d:data=8'h00;
14'h2b7e:data=8'h00;
14'h2b7f:data=8'h00;
14'h3300:data=8'h00;
14'h3301:data=8'h00;
14'h3302:data=8'h00;
14'h3303:data=8'h00;
14'h3304:data=8'h00;
14'h3305:data=8'h00;
14'h3306:data=8'h00;
14'h3307:data=8'h00;
14'h3308:data=8'h00;
14'h3309:data=8'h00;
14'h330a:data=8'h00;
14'h330b:data=8'h00;
14'h330c:data=8'h00;
14'h330d:data=8'h00;
14'h330e:data=8'h00;
14'h330f:data=8'h00;
14'h3310:data=8'h00;
14'h3311:data=8'h00;
14'h3312:data=8'h00;
14'h3313:data=8'h00;
14'h3314:data=8'h00;
14'h3315:data=8'h00;
14'h3316:data=8'h00;
14'h3317:data=8'h00;
14'h3318:data=8'h00;
14'h3319:data=8'h00;
14'h331a:data=8'h00;
14'h331b:data=8'h00;
14'h331c:data=8'h00;
14'h331d:data=8'h00;
14'h331e:data=8'h00;
14'h331f:data=8'h00;
14'h3320:data=8'h00;
14'h3321:data=8'h00;
14'h3322:data=8'h00;
14'h3323:data=8'h00;
14'h3324:data=8'h00;
14'h3325:data=8'h00;
14'h3326:data=8'h00;
14'h3327:data=8'h00;
14'h3328:data=8'h00;
14'h3329:data=8'h00;
14'h332a:data=8'h00;
14'h332b:data=8'h00;
14'h332c:data=8'h00;
14'h332d:data=8'h00;
14'h332e:data=8'hFC;
14'h332f:data=8'hFF;
14'h3330:data=8'hFF;
14'h3331:data=8'hFF;
14'h3332:data=8'hFE;
14'h3333:data=8'hFE;
14'h3334:data=8'hFE;
14'h3335:data=8'hFC;
14'h3336:data=8'hFC;
14'h3337:data=8'hFE;
14'h3338:data=8'hFE;
14'h3339:data=8'hFF;
14'h333a:data=8'hFF;
14'h333b:data=8'hFF;
14'h333c:data=8'hFF;
14'h333d:data=8'hFF;
14'h333e:data=8'h7F;
14'h333f:data=8'h7F;
14'h3340:data=8'h3F;
14'h3341:data=8'h1F;
14'h3342:data=8'h07;
14'h3343:data=8'h01;
14'h3344:data=8'h00;
14'h3345:data=8'h00;
14'h3346:data=8'h00;
14'h3347:data=8'h00;
14'h3348:data=8'h00;
14'h3349:data=8'h00;
14'h334a:data=8'h00;
14'h334b:data=8'h00;
14'h334c:data=8'h00;
14'h334d:data=8'h00;
14'h334e:data=8'h00;
14'h334f:data=8'h00;
14'h3350:data=8'h00;
14'h3351:data=8'h00;
14'h3352:data=8'h00;
14'h3353:data=8'h00;
14'h3354:data=8'h00;
14'h3355:data=8'h00;
14'h3356:data=8'h00;
14'h3357:data=8'h00;
14'h3358:data=8'h00;
14'h3359:data=8'h00;
14'h335a:data=8'h00;
14'h335b:data=8'h00;
14'h335c:data=8'h00;
14'h335d:data=8'h00;
14'h335e:data=8'h00;
14'h335f:data=8'h00;
14'h3360:data=8'h00;
14'h3361:data=8'h00;
14'h3362:data=8'h00;
14'h3363:data=8'h00;
14'h3364:data=8'h00;
14'h3365:data=8'h00;
14'h3366:data=8'h00;
14'h3367:data=8'h00;
14'h3368:data=8'h00;
14'h3369:data=8'h00;
14'h336a:data=8'h00;
14'h336b:data=8'h00;
14'h336c:data=8'h00;
14'h336d:data=8'h00;
14'h336e:data=8'h00;
14'h336f:data=8'h00;
14'h3370:data=8'h00;
14'h3371:data=8'h00;
14'h3372:data=8'h00;
14'h3373:data=8'h00;
14'h3374:data=8'h00;
14'h3375:data=8'h00;
14'h3376:data=8'h00;
14'h3377:data=8'h00;
14'h3378:data=8'h00;
14'h3379:data=8'h00;
14'h337a:data=8'h00;
14'h337b:data=8'h00;
14'h337c:data=8'h00;
14'h337d:data=8'h00;
14'h337e:data=8'h00;
14'h337f:data=8'h00;
14'h3b00:data=8'h00;
14'h3b01:data=8'h00;
14'h3b02:data=8'h00;
14'h3b03:data=8'h00;
14'h3b04:data=8'h00;
14'h3b05:data=8'h00;
14'h3b06:data=8'h00;
14'h3b07:data=8'h00;
14'h3b08:data=8'h00;
14'h3b09:data=8'h00;
14'h3b0a:data=8'h00;
14'h3b0b:data=8'h00;
14'h3b0c:data=8'h00;
14'h3b0d:data=8'h00;
14'h3b0e:data=8'h00;
14'h3b0f:data=8'h00;
14'h3b10:data=8'h00;
14'h3b11:data=8'h00;
14'h3b12:data=8'h00;
14'h3b13:data=8'h00;
14'h3b14:data=8'h00;
14'h3b15:data=8'h00;
14'h3b16:data=8'h00;
14'h3b17:data=8'h00;
14'h3b18:data=8'h00;
14'h3b19:data=8'h00;
14'h3b1a:data=8'h00;
14'h3b1b:data=8'h00;
14'h3b1c:data=8'h00;
14'h3b1d:data=8'h00;
14'h3b1e:data=8'h00;
14'h3b1f:data=8'h00;
14'h3b20:data=8'h00;
14'h3b21:data=8'h00;
14'h3b22:data=8'h00;
14'h3b23:data=8'h00;
14'h3b24:data=8'h00;
14'h3b25:data=8'h00;
14'h3b26:data=8'h00;
14'h3b27:data=8'h00;
14'h3b28:data=8'h00;
14'h3b29:data=8'h00;
14'h3b2a:data=8'h00;
14'h3b2b:data=8'h00;
14'h3b2c:data=8'h00;
14'h3b2d:data=8'h00;
14'h3b2e:data=8'h00;
14'h3b2f:data=8'h00;
14'h3b30:data=8'h01;
14'h3b31:data=8'h01;
14'h3b32:data=8'h01;
14'h3b33:data=8'h01;
14'h3b34:data=8'h01;
14'h3b35:data=8'h01;
14'h3b36:data=8'h01;
14'h3b37:data=8'h01;
14'h3b38:data=8'h01;
14'h3b39:data=8'h01;
14'h3b3a:data=8'h01;
14'h3b3b:data=8'h01;
14'h3b3c:data=8'h00;
14'h3b3d:data=8'h00;
14'h3b3e:data=8'h00;
14'h3b3f:data=8'h00;
14'h3b40:data=8'h00;
14'h3b41:data=8'h00;
14'h3b42:data=8'h00;
14'h3b43:data=8'h00;
14'h3b44:data=8'h00;
14'h3b45:data=8'h00;
14'h3b46:data=8'h00;
14'h3b47:data=8'h00;
14'h3b48:data=8'h00;
14'h3b49:data=8'h00;
14'h3b4a:data=8'h00;
14'h3b4b:data=8'h00;
14'h3b4c:data=8'h00;
14'h3b4d:data=8'h00;
14'h3b4e:data=8'h00;
14'h3b4f:data=8'h00;
14'h3b50:data=8'h00;
14'h3b51:data=8'h00;
14'h3b52:data=8'h00;
14'h3b53:data=8'h00;
14'h3b54:data=8'h00;
14'h3b55:data=8'h00;
14'h3b56:data=8'h00;
14'h3b57:data=8'h00;
14'h3b58:data=8'h00;
14'h3b59:data=8'h00;
14'h3b5a:data=8'h00;
14'h3b5b:data=8'h00;
14'h3b5c:data=8'h00;
14'h3b5d:data=8'h00;
14'h3b5e:data=8'h00;
14'h3b5f:data=8'h00;
14'h3b60:data=8'h00;
14'h3b61:data=8'h00;
14'h3b62:data=8'h00;
14'h3b63:data=8'h00;
14'h3b64:data=8'h00;
14'h3b65:data=8'h00;
14'h3b66:data=8'h00;
14'h3b67:data=8'h00;
14'h3b68:data=8'h00;
14'h3b69:data=8'h00;
14'h3b6a:data=8'h00;
14'h3b6b:data=8'h00;
14'h3b6c:data=8'h00;
14'h3b6d:data=8'h00;
14'h3b6e:data=8'h00;
14'h3b6f:data=8'h00;
14'h3b70:data=8'h00;
14'h3b71:data=8'h00;
14'h3b72:data=8'h00;
14'h3b73:data=8'h00;
14'h3b74:data=8'h00;
14'h3b75:data=8'h00;
14'h3b76:data=8'h00;
14'h3b77:data=8'h00;
14'h3b78:data=8'h00;
14'h3b79:data=8'h00;
14'h3b7a:data=8'h00;
14'h3b7b:data=8'h00;
14'h3b7c:data=8'h00;
14'h3b7d:data=8'h00;
14'h3b7e:data=8'h00;
14'h3b7f:data=8'h00;
////////////////////////////////////////////////////////////////////////////////////////PIC5 Info
14'h0400:data=8'h00;
14'h0401:data=8'h00;
14'h0402:data=8'h00;
14'h0403:data=8'h00;
14'h0404:data=8'h00;
14'h0405:data=8'h00;
14'h0406:data=8'h00;
14'h0407:data=8'h00;
14'h0408:data=8'h00;
14'h0409:data=8'h00;
14'h040a:data=8'h00;
14'h040b:data=8'h00;
14'h040c:data=8'h00;
14'h040d:data=8'h00;
14'h040e:data=8'h00;
14'h040f:data=8'h00;
14'h0410:data=8'h00;
14'h0411:data=8'h00;
14'h0412:data=8'h00;
14'h0413:data=8'h00;
14'h0414:data=8'h00;
14'h0415:data=8'h00;
14'h0416:data=8'h00;
14'h0417:data=8'h00;
14'h0418:data=8'h00;
14'h0419:data=8'h00;
14'h041a:data=8'h00;
14'h041b:data=8'h00;
14'h041c:data=8'h00;
14'h041d:data=8'h00;
14'h041e:data=8'h00;
14'h041f:data=8'h00;
14'h0420:data=8'h00;
14'h0421:data=8'h00;
14'h0422:data=8'h00;
14'h0423:data=8'h00;
14'h0424:data=8'h00;
14'h0425:data=8'h00;
14'h0426:data=8'h00;
14'h0427:data=8'h00;
14'h0428:data=8'h00;
14'h0429:data=8'h00;
14'h042a:data=8'h00;
14'h042b:data=8'h00;
14'h042c:data=8'h00;
14'h042d:data=8'h00;
14'h042e:data=8'h00;
14'h042f:data=8'h00;
14'h0430:data=8'h00;
14'h0431:data=8'h00;
14'h0432:data=8'h00;
14'h0433:data=8'h00;
14'h0434:data=8'h00;
14'h0435:data=8'h00;
14'h0436:data=8'h00;
14'h0437:data=8'h00;
14'h0438:data=8'h00;
14'h0439:data=8'h00;
14'h043a:data=8'h00;
14'h043b:data=8'h00;
14'h043c:data=8'h00;
14'h043d:data=8'h00;
14'h043e:data=8'h00;
14'h043f:data=8'h00;
14'h0440:data=8'h00;
14'h0441:data=8'h00;
14'h0442:data=8'h00;
14'h0443:data=8'h00;
14'h0444:data=8'h00;
14'h0445:data=8'h00;
14'h0446:data=8'h00;
14'h0447:data=8'h00;
14'h0448:data=8'h00;
14'h0449:data=8'h00;
14'h044a:data=8'h00;
14'h044b:data=8'h00;
14'h044c:data=8'h00;
14'h044d:data=8'h00;
14'h044e:data=8'h00;
14'h044f:data=8'h00;
14'h0450:data=8'h00;
14'h0451:data=8'h00;
14'h0452:data=8'h00;
14'h0453:data=8'h00;
14'h0454:data=8'h00;
14'h0455:data=8'h00;
14'h0456:data=8'h00;
14'h0457:data=8'h00;
14'h0458:data=8'h00;
14'h0459:data=8'h00;
14'h045a:data=8'h00;
14'h045b:data=8'h00;
14'h045c:data=8'h00;
14'h045d:data=8'h00;
14'h045e:data=8'h00;
14'h045f:data=8'h00;
14'h0460:data=8'h00;
14'h0461:data=8'h00;
14'h0462:data=8'h00;
14'h0463:data=8'h00;
14'h0464:data=8'h00;
14'h0465:data=8'h00;
14'h0466:data=8'h00;
14'h0467:data=8'h00;
14'h0468:data=8'h00;
14'h0469:data=8'h00;
14'h046a:data=8'h00;
14'h046b:data=8'h00;
14'h046c:data=8'h00;
14'h046d:data=8'h00;
14'h046e:data=8'h00;
14'h046f:data=8'h00;
14'h0470:data=8'h00;
14'h0471:data=8'h00;
14'h0472:data=8'h00;
14'h0473:data=8'h00;
14'h0474:data=8'h00;
14'h0475:data=8'h00;
14'h0476:data=8'h00;
14'h0477:data=8'h00;
14'h0478:data=8'h00;
14'h0479:data=8'h00;
14'h047a:data=8'h00;
14'h047b:data=8'h00;
14'h047c:data=8'h00;
14'h047d:data=8'h00;
14'h047e:data=8'h00;
14'h047f:data=8'h00;
14'h0c00:data=8'h00;
14'h0c01:data=8'h00;
14'h0c02:data=8'h00;
14'h0c03:data=8'h00;
14'h0c04:data=8'h00;
14'h0c05:data=8'h00;
14'h0c06:data=8'h00;
14'h0c07:data=8'h00;
14'h0c08:data=8'h00;
14'h0c09:data=8'h00;
14'h0c0a:data=8'h00;
14'h0c0b:data=8'h00;
14'h0c0c:data=8'h00;
14'h0c0d:data=8'h00;
14'h0c0e:data=8'h00;
14'h0c0f:data=8'h00;
14'h0c10:data=8'h00;
14'h0c11:data=8'h00;
14'h0c12:data=8'h00;
14'h0c13:data=8'h00;
14'h0c14:data=8'h00;
14'h0c15:data=8'h00;
14'h0c16:data=8'h00;
14'h0c17:data=8'h00;
14'h0c18:data=8'h00;
14'h0c19:data=8'h00;
14'h0c1a:data=8'h00;
14'h0c1b:data=8'h00;
14'h0c1c:data=8'h00;
14'h0c1d:data=8'h00;
14'h0c1e:data=8'h00;
14'h0c1f:data=8'h00;
14'h0c20:data=8'h00;
14'h0c21:data=8'h00;
14'h0c22:data=8'h00;
14'h0c23:data=8'h00;
14'h0c24:data=8'h00;
14'h0c25:data=8'h00;
14'h0c26:data=8'h00;
14'h0c27:data=8'h00;
14'h0c28:data=8'h00;
14'h0c29:data=8'h00;
14'h0c2a:data=8'h00;
14'h0c2b:data=8'h00;
14'h0c2c:data=8'h00;
14'h0c2d:data=8'h00;
14'h0c2e:data=8'h00;
14'h0c2f:data=8'h00;
14'h0c30:data=8'h00;
14'h0c31:data=8'h00;
14'h0c32:data=8'h00;
14'h0c33:data=8'h00;
14'h0c34:data=8'h00;
14'h0c35:data=8'h00;
14'h0c36:data=8'h00;
14'h0c37:data=8'h00;
14'h0c38:data=8'h00;
14'h0c39:data=8'h00;
14'h0c3a:data=8'h00;
14'h0c3b:data=8'h00;
14'h0c3c:data=8'h00;
14'h0c3d:data=8'h00;
14'h0c3e:data=8'h00;
14'h0c3f:data=8'h00;
14'h0c40:data=8'h00;
14'h0c41:data=8'h00;
14'h0c42:data=8'h00;
14'h0c43:data=8'h00;
14'h0c44:data=8'h00;
14'h0c45:data=8'h80;
14'h0c46:data=8'h80;
14'h0c47:data=8'hC0;
14'h0c48:data=8'hC0;
14'h0c49:data=8'hC0;
14'h0c4a:data=8'hC0;
14'h0c4b:data=8'hC0;
14'h0c4c:data=8'hC0;
14'h0c4d:data=8'hC0;
14'h0c4e:data=8'hC0;
14'h0c4f:data=8'hC0;
14'h0c50:data=8'hC0;
14'h0c51:data=8'h00;
14'h0c52:data=8'h00;
14'h0c53:data=8'h00;
14'h0c54:data=8'h00;
14'h0c55:data=8'h00;
14'h0c56:data=8'h00;
14'h0c57:data=8'h00;
14'h0c58:data=8'h00;
14'h0c59:data=8'h00;
14'h0c5a:data=8'h00;
14'h0c5b:data=8'h00;
14'h0c5c:data=8'h00;
14'h0c5d:data=8'h00;
14'h0c5e:data=8'h00;
14'h0c5f:data=8'h00;
14'h0c60:data=8'h00;
14'h0c61:data=8'h00;
14'h0c62:data=8'h00;
14'h0c63:data=8'h00;
14'h0c64:data=8'h00;
14'h0c65:data=8'h00;
14'h0c66:data=8'h00;
14'h0c67:data=8'h00;
14'h0c68:data=8'h00;
14'h0c69:data=8'h00;
14'h0c6a:data=8'h00;
14'h0c6b:data=8'h00;
14'h0c6c:data=8'h00;
14'h0c6d:data=8'h00;
14'h0c6e:data=8'h00;
14'h0c6f:data=8'h00;
14'h0c70:data=8'h00;
14'h0c71:data=8'h00;
14'h0c72:data=8'h00;
14'h0c73:data=8'h00;
14'h0c74:data=8'h00;
14'h0c75:data=8'h00;
14'h0c76:data=8'h00;
14'h0c77:data=8'h00;
14'h0c78:data=8'h00;
14'h0c79:data=8'h00;
14'h0c7a:data=8'h00;
14'h0c7b:data=8'h00;
14'h0c7c:data=8'h00;
14'h0c7d:data=8'h00;
14'h0c7e:data=8'h00;
14'h0c7f:data=8'h00;
14'h1400:data=8'h00;
14'h1401:data=8'h00;
14'h1402:data=8'h00;
14'h1403:data=8'h00;
14'h1404:data=8'h00;
14'h1405:data=8'h00;
14'h1406:data=8'h00;
14'h1407:data=8'h00;
14'h1408:data=8'h00;
14'h1409:data=8'h00;
14'h140a:data=8'h00;
14'h140b:data=8'h00;
14'h140c:data=8'h00;
14'h140d:data=8'h00;
14'h140e:data=8'h00;
14'h140f:data=8'h00;
14'h1410:data=8'h00;
14'h1411:data=8'h00;
14'h1412:data=8'h00;
14'h1413:data=8'h00;
14'h1414:data=8'h00;
14'h1415:data=8'h00;
14'h1416:data=8'h00;
14'h1417:data=8'h00;
14'h1418:data=8'h00;
14'h1419:data=8'h00;
14'h141a:data=8'h00;
14'h141b:data=8'hC0;
14'h141c:data=8'hFC;
14'h141d:data=8'hFF;
14'h141e:data=8'hFF;
14'h141f:data=8'hFF;
14'h1420:data=8'hFF;
14'h1421:data=8'hFF;
14'h1422:data=8'hFF;
14'h1423:data=8'hFF;
14'h1424:data=8'h3F;
14'h1425:data=8'h00;
14'h1426:data=8'h00;
14'h1427:data=8'h00;
14'h1428:data=8'h00;
14'h1429:data=8'h00;
14'h142a:data=8'h00;
14'h142b:data=8'h00;
14'h142c:data=8'h00;
14'h142d:data=8'h00;
14'h142e:data=8'h00;
14'h142f:data=8'h00;
14'h1430:data=8'h00;
14'h1431:data=8'h00;
14'h1432:data=8'h00;
14'h1433:data=8'h00;
14'h1434:data=8'h00;
14'h1435:data=8'h00;
14'h1436:data=8'h00;
14'h1437:data=8'h00;
14'h1438:data=8'h00;
14'h1439:data=8'h00;
14'h143a:data=8'h00;
14'h143b:data=8'h00;
14'h143c:data=8'h00;
14'h143d:data=8'h00;
14'h143e:data=8'h00;
14'h143f:data=8'h00;
14'h1440:data=8'h00;
14'h1441:data=8'h80;
14'h1442:data=8'hF8;
14'h1443:data=8'hFE;
14'h1444:data=8'hFF;
14'h1445:data=8'hFF;
14'h1446:data=8'hFF;
14'h1447:data=8'hFF;
14'h1448:data=8'hFF;
14'h1449:data=8'hFF;
14'h144a:data=8'h7F;
14'h144b:data=8'h3F;
14'h144c:data=8'h1F;
14'h144d:data=8'h3F;
14'h144e:data=8'h3F;
14'h144f:data=8'h3F;
14'h1450:data=8'h0F;
14'h1451:data=8'h00;
14'h1452:data=8'h00;
14'h1453:data=8'h00;
14'h1454:data=8'h00;
14'h1455:data=8'h00;
14'h1456:data=8'h00;
14'h1457:data=8'h00;
14'h1458:data=8'h00;
14'h1459:data=8'h00;
14'h145a:data=8'h00;
14'h145b:data=8'h00;
14'h145c:data=8'h00;
14'h145d:data=8'h00;
14'h145e:data=8'h00;
14'h145f:data=8'h00;
14'h1460:data=8'h00;
14'h1461:data=8'h00;
14'h1462:data=8'h00;
14'h1463:data=8'h00;
14'h1464:data=8'h00;
14'h1465:data=8'h00;
14'h1466:data=8'h00;
14'h1467:data=8'h00;
14'h1468:data=8'h00;
14'h1469:data=8'h00;
14'h146a:data=8'h00;
14'h146b:data=8'h00;
14'h146c:data=8'h00;
14'h146d:data=8'h00;
14'h146e:data=8'h00;
14'h146f:data=8'h00;
14'h1470:data=8'h00;
14'h1471:data=8'h00;
14'h1472:data=8'h00;
14'h1473:data=8'h00;
14'h1474:data=8'h00;
14'h1475:data=8'h00;
14'h1476:data=8'h00;
14'h1477:data=8'h00;
14'h1478:data=8'h00;
14'h1479:data=8'h00;
14'h147a:data=8'h00;
14'h147b:data=8'h00;
14'h147c:data=8'h00;
14'h147d:data=8'h00;
14'h147e:data=8'h00;
14'h147f:data=8'h00;
14'h1c00:data=8'h00;
14'h1c01:data=8'h00;
14'h1c02:data=8'h00;
14'h1c03:data=8'h00;
14'h1c04:data=8'h00;
14'h1c05:data=8'h00;
14'h1c06:data=8'h00;
14'h1c07:data=8'h00;
14'h1c08:data=8'h00;
14'h1c09:data=8'h00;
14'h1c0a:data=8'h00;
14'h1c0b:data=8'h00;
14'h1c0c:data=8'h00;
14'h1c0d:data=8'h00;
14'h1c0e:data=8'h00;
14'h1c0f:data=8'h00;
14'h1c10:data=8'h00;
14'h1c11:data=8'h00;
14'h1c12:data=8'h00;
14'h1c13:data=8'h00;
14'h1c14:data=8'h00;
14'h1c15:data=8'h00;
14'h1c16:data=8'h00;
14'h1c17:data=8'h00;
14'h1c18:data=8'h00;
14'h1c19:data=8'h00;
14'h1c1a:data=8'hF8;
14'h1c1b:data=8'hFF;
14'h1c1c:data=8'hFF;
14'h1c1d:data=8'hFF;
14'h1c1e:data=8'hFF;
14'h1c1f:data=8'hFF;
14'h1c20:data=8'hFF;
14'h1c21:data=8'hFF;
14'h1c22:data=8'hFF;
14'h1c23:data=8'h07;
14'h1c24:data=8'h00;
14'h1c25:data=8'h00;
14'h1c26:data=8'hC0;
14'h1c27:data=8'hFF;
14'h1c28:data=8'hFF;
14'h1c29:data=8'hFF;
14'h1c2a:data=8'hFF;
14'h1c2b:data=8'hFF;
14'h1c2c:data=8'hFF;
14'h1c2d:data=8'hFF;
14'h1c2e:data=8'hFF;
14'h1c2f:data=8'hFF;
14'h1c30:data=8'hFE;
14'h1c31:data=8'hFF;
14'h1c32:data=8'hFF;
14'h1c33:data=8'hFF;
14'h1c34:data=8'hFF;
14'h1c35:data=8'hFF;
14'h1c36:data=8'hFF;
14'h1c37:data=8'hFF;
14'h1c38:data=8'hFF;
14'h1c39:data=8'hFF;
14'h1c3a:data=8'hFC;
14'h1c3b:data=8'h00;
14'h1c3c:data=8'h00;
14'h1c3d:data=8'h7E;
14'h1c3e:data=8'h7F;
14'h1c3f:data=8'h7F;
14'h1c40:data=8'hFF;
14'h1c41:data=8'hFF;
14'h1c42:data=8'hFF;
14'h1c43:data=8'hFF;
14'h1c44:data=8'hFF;
14'h1c45:data=8'hFF;
14'h1c46:data=8'hFF;
14'h1c47:data=8'hFF;
14'h1c48:data=8'hFF;
14'h1c49:data=8'h7F;
14'h1c4a:data=8'h7F;
14'h1c4b:data=8'h7F;
14'h1c4c:data=8'h7F;
14'h1c4d:data=8'hFF;
14'h1c4e:data=8'hE0;
14'h1c4f:data=8'hF8;
14'h1c50:data=8'hFC;
14'h1c51:data=8'hFC;
14'h1c52:data=8'hFE;
14'h1c53:data=8'hFE;
14'h1c54:data=8'hFF;
14'h1c55:data=8'hFF;
14'h1c56:data=8'hFF;
14'h1c57:data=8'hFF;
14'h1c58:data=8'hFF;
14'h1c59:data=8'h7F;
14'h1c5a:data=8'hFF;
14'h1c5b:data=8'hFF;
14'h1c5c:data=8'hFF;
14'h1c5d:data=8'hFF;
14'h1c5e:data=8'hFF;
14'h1c5f:data=8'hFE;
14'h1c60:data=8'hFE;
14'h1c61:data=8'hFC;
14'h1c62:data=8'hF0;
14'h1c63:data=8'h00;
14'h1c64:data=8'h00;
14'h1c65:data=8'h00;
14'h1c66:data=8'h00;
14'h1c67:data=8'h00;
14'h1c68:data=8'h00;
14'h1c69:data=8'h00;
14'h1c6a:data=8'h00;
14'h1c6b:data=8'h00;
14'h1c6c:data=8'h00;
14'h1c6d:data=8'h00;
14'h1c6e:data=8'h00;
14'h1c6f:data=8'h00;
14'h1c70:data=8'h00;
14'h1c71:data=8'h00;
14'h1c72:data=8'h00;
14'h1c73:data=8'h00;
14'h1c74:data=8'h00;
14'h1c75:data=8'h00;
14'h1c76:data=8'h00;
14'h1c77:data=8'h00;
14'h1c78:data=8'h00;
14'h1c79:data=8'h00;
14'h1c7a:data=8'h00;
14'h1c7b:data=8'h00;
14'h1c7c:data=8'h00;
14'h1c7d:data=8'h00;
14'h1c7e:data=8'h00;
14'h1c7f:data=8'h00;
14'h2400:data=8'h00;
14'h2401:data=8'h00;
14'h2402:data=8'h00;
14'h2403:data=8'h00;
14'h2404:data=8'h00;
14'h2405:data=8'h00;
14'h2406:data=8'h00;
14'h2407:data=8'h00;
14'h2408:data=8'h00;
14'h2409:data=8'h00;
14'h240a:data=8'h00;
14'h240b:data=8'h00;
14'h240c:data=8'h00;
14'h240d:data=8'h00;
14'h240e:data=8'h00;
14'h240f:data=8'h00;
14'h2410:data=8'h00;
14'h2411:data=8'h00;
14'h2412:data=8'h00;
14'h2413:data=8'h00;
14'h2414:data=8'h00;
14'h2415:data=8'h00;
14'h2416:data=8'h00;
14'h2417:data=8'h00;
14'h2418:data=8'hE0;
14'h2419:data=8'hFF;
14'h241a:data=8'hFF;
14'h241b:data=8'hFF;
14'h241c:data=8'hFF;
14'h241d:data=8'hFF;
14'h241e:data=8'hFF;
14'h241f:data=8'hFF;
14'h2420:data=8'hFF;
14'h2421:data=8'h0F;
14'h2422:data=8'h00;
14'h2423:data=8'h00;
14'h2424:data=8'h80;
14'h2425:data=8'hF8;
14'h2426:data=8'hFF;
14'h2427:data=8'hFF;
14'h2428:data=8'hFF;
14'h2429:data=8'hFF;
14'h242a:data=8'hFF;
14'h242b:data=8'hFF;
14'h242c:data=8'hFF;
14'h242d:data=8'h7F;
14'h242e:data=8'h0F;
14'h242f:data=8'h03;
14'h2430:data=8'h01;
14'h2431:data=8'h00;
14'h2432:data=8'hE0;
14'h2433:data=8'hFF;
14'h2434:data=8'hFF;
14'h2435:data=8'hFF;
14'h2436:data=8'hFF;
14'h2437:data=8'hFF;
14'h2438:data=8'hFF;
14'h2439:data=8'hFF;
14'h243a:data=8'h0F;
14'h243b:data=8'h00;
14'h243c:data=8'h00;
14'h243d:data=8'h00;
14'h243e:data=8'hE0;
14'h243f:data=8'hFF;
14'h2440:data=8'hFF;
14'h2441:data=8'hFF;
14'h2442:data=8'hFF;
14'h2443:data=8'hFF;
14'h2444:data=8'hFF;
14'h2445:data=8'hFF;
14'h2446:data=8'hFF;
14'h2447:data=8'h0F;
14'h2448:data=8'h00;
14'h2449:data=8'h00;
14'h244a:data=8'h00;
14'h244b:data=8'h00;
14'h244c:data=8'hFE;
14'h244d:data=8'hFF;
14'h244e:data=8'hFF;
14'h244f:data=8'hFF;
14'h2450:data=8'hFF;
14'h2451:data=8'hFF;
14'h2452:data=8'hFF;
14'h2453:data=8'hFF;
14'h2454:data=8'hFF;
14'h2455:data=8'h03;
14'h2456:data=8'h01;
14'h2457:data=8'h00;
14'h2458:data=8'h00;
14'h2459:data=8'h80;
14'h245a:data=8'hE0;
14'h245b:data=8'hFF;
14'h245c:data=8'hFF;
14'h245d:data=8'hFF;
14'h245e:data=8'hFF;
14'h245f:data=8'hFF;
14'h2460:data=8'hFF;
14'h2461:data=8'hFF;
14'h2462:data=8'hFF;
14'h2463:data=8'h0F;
14'h2464:data=8'h00;
14'h2465:data=8'h00;
14'h2466:data=8'h00;
14'h2467:data=8'h00;
14'h2468:data=8'h00;
14'h2469:data=8'h00;
14'h246a:data=8'h00;
14'h246b:data=8'h00;
14'h246c:data=8'h00;
14'h246d:data=8'h00;
14'h246e:data=8'h00;
14'h246f:data=8'h00;
14'h2470:data=8'h00;
14'h2471:data=8'h00;
14'h2472:data=8'h00;
14'h2473:data=8'h00;
14'h2474:data=8'h00;
14'h2475:data=8'h00;
14'h2476:data=8'h00;
14'h2477:data=8'h00;
14'h2478:data=8'h00;
14'h2479:data=8'h00;
14'h247a:data=8'h00;
14'h247b:data=8'h00;
14'h247c:data=8'h00;
14'h247d:data=8'h00;
14'h247e:data=8'h00;
14'h247f:data=8'h00;
14'h2c00:data=8'h00;
14'h2c01:data=8'h00;
14'h2c02:data=8'h00;
14'h2c03:data=8'h00;
14'h2c04:data=8'h00;
14'h2c05:data=8'h00;
14'h2c06:data=8'h00;
14'h2c07:data=8'h00;
14'h2c08:data=8'h00;
14'h2c09:data=8'h00;
14'h2c0a:data=8'h00;
14'h2c0b:data=8'h00;
14'h2c0c:data=8'h00;
14'h2c0d:data=8'h00;
14'h2c0e:data=8'h00;
14'h2c0f:data=8'h00;
14'h2c10:data=8'h00;
14'h2c11:data=8'h00;
14'h2c12:data=8'h00;
14'h2c13:data=8'h00;
14'h2c14:data=8'h00;
14'h2c15:data=8'h00;
14'h2c16:data=8'h00;
14'h2c17:data=8'h00;
14'h2c18:data=8'h7F;
14'h2c19:data=8'h7F;
14'h2c1a:data=8'h7F;
14'h2c1b:data=8'h7F;
14'h2c1c:data=8'h7F;
14'h2c1d:data=8'h7F;
14'h2c1e:data=8'h7F;
14'h2c1f:data=8'h1F;
14'h2c20:data=8'h01;
14'h2c21:data=8'h00;
14'h2c22:data=8'h00;
14'h2c23:data=8'h70;
14'h2c24:data=8'h7F;
14'h2c25:data=8'h7F;
14'h2c26:data=8'h7F;
14'h2c27:data=8'h7F;
14'h2c28:data=8'h7F;
14'h2c29:data=8'h7F;
14'h2c2a:data=8'h7F;
14'h2c2b:data=8'h7F;
14'h2c2c:data=8'h07;
14'h2c2d:data=8'h00;
14'h2c2e:data=8'h00;
14'h2c2f:data=8'h00;
14'h2c30:data=8'h00;
14'h2c31:data=8'h7C;
14'h2c32:data=8'h7F;
14'h2c33:data=8'h7F;
14'h2c34:data=8'h7F;
14'h2c35:data=8'h7F;
14'h2c36:data=8'h7F;
14'h2c37:data=8'h7F;
14'h2c38:data=8'h7F;
14'h2c39:data=8'h1F;
14'h2c3a:data=8'h00;
14'h2c3b:data=8'h00;
14'h2c3c:data=8'h80;
14'h2c3d:data=8'hFC;
14'h2c3e:data=8'hFF;
14'h2c3f:data=8'hFF;
14'h2c40:data=8'hFF;
14'h2c41:data=8'hFF;
14'h2c42:data=8'hFF;
14'h2c43:data=8'hFF;
14'h2c44:data=8'hFF;
14'h2c45:data=8'h1F;
14'h2c46:data=8'h01;
14'h2c47:data=8'h00;
14'h2c48:data=8'h00;
14'h2c49:data=8'h00;
14'h2c4a:data=8'h00;
14'h2c4b:data=8'h00;
14'h2c4c:data=8'h01;
14'h2c4d:data=8'h0F;
14'h2c4e:data=8'h1F;
14'h2c4f:data=8'h3F;
14'h2c50:data=8'h3F;
14'h2c51:data=8'h7F;
14'h2c52:data=8'h7F;
14'h2c53:data=8'h7F;
14'h2c54:data=8'h7F;
14'h2c55:data=8'h7F;
14'h2c56:data=8'h7F;
14'h2c57:data=8'h7F;
14'h2c58:data=8'h7F;
14'h2c59:data=8'h7F;
14'h2c5a:data=8'h7F;
14'h2c5b:data=8'h7F;
14'h2c5c:data=8'h3F;
14'h2c5d:data=8'h3F;
14'h2c5e:data=8'h1F;
14'h2c5f:data=8'h0F;
14'h2c60:data=8'h07;
14'h2c61:data=8'h03;
14'h2c62:data=8'h00;
14'h2c63:data=8'h00;
14'h2c64:data=8'h00;
14'h2c65:data=8'h00;
14'h2c66:data=8'h00;
14'h2c67:data=8'h00;
14'h2c68:data=8'h00;
14'h2c69:data=8'h00;
14'h2c6a:data=8'h00;
14'h2c6b:data=8'h00;
14'h2c6c:data=8'h00;
14'h2c6d:data=8'h00;
14'h2c6e:data=8'h00;
14'h2c6f:data=8'h00;
14'h2c70:data=8'h00;
14'h2c71:data=8'h00;
14'h2c72:data=8'h00;
14'h2c73:data=8'h00;
14'h2c74:data=8'h00;
14'h2c75:data=8'h00;
14'h2c76:data=8'h00;
14'h2c77:data=8'h00;
14'h2c78:data=8'h00;
14'h2c79:data=8'h00;
14'h2c7a:data=8'h00;
14'h2c7b:data=8'h00;
14'h2c7c:data=8'h00;
14'h2c7d:data=8'h00;
14'h2c7e:data=8'h00;
14'h2c7f:data=8'h00;
14'h3400:data=8'h00;
14'h3401:data=8'h00;
14'h3402:data=8'h00;
14'h3403:data=8'h00;
14'h3404:data=8'h00;
14'h3405:data=8'h00;
14'h3406:data=8'h00;
14'h3407:data=8'h00;
14'h3408:data=8'h00;
14'h3409:data=8'h00;
14'h340a:data=8'h00;
14'h340b:data=8'h00;
14'h340c:data=8'h00;
14'h340d:data=8'h00;
14'h340e:data=8'h00;
14'h340f:data=8'h00;
14'h3410:data=8'h00;
14'h3411:data=8'h00;
14'h3412:data=8'h00;
14'h3413:data=8'h00;
14'h3414:data=8'h00;
14'h3415:data=8'h00;
14'h3416:data=8'h00;
14'h3417:data=8'h00;
14'h3418:data=8'h00;
14'h3419:data=8'h00;
14'h341a:data=8'h00;
14'h341b:data=8'h00;
14'h341c:data=8'h00;
14'h341d:data=8'h00;
14'h341e:data=8'h00;
14'h341f:data=8'h00;
14'h3420:data=8'h00;
14'h3421:data=8'h00;
14'h3422:data=8'h00;
14'h3423:data=8'h00;
14'h3424:data=8'h00;
14'h3425:data=8'h00;
14'h3426:data=8'h00;
14'h3427:data=8'h00;
14'h3428:data=8'h00;
14'h3429:data=8'h00;
14'h342a:data=8'h00;
14'h342b:data=8'h00;
14'h342c:data=8'h00;
14'h342d:data=8'h00;
14'h342e:data=8'h00;
14'h342f:data=8'h00;
14'h3430:data=8'h00;
14'h3431:data=8'h00;
14'h3432:data=8'h00;
14'h3433:data=8'h00;
14'h3434:data=8'h00;
14'h3435:data=8'h00;
14'h3436:data=8'h00;
14'h3437:data=8'h00;
14'h3438:data=8'h00;
14'h3439:data=8'h00;
14'h343a:data=8'h00;
14'h343b:data=8'h38;
14'h343c:data=8'h3F;
14'h343d:data=8'h3F;
14'h343e:data=8'h3F;
14'h343f:data=8'h3F;
14'h3440:data=8'h3F;
14'h3441:data=8'h3F;
14'h3442:data=8'h3F;
14'h3443:data=8'h3F;
14'h3444:data=8'h03;
14'h3445:data=8'h00;
14'h3446:data=8'h00;
14'h3447:data=8'h00;
14'h3448:data=8'h00;
14'h3449:data=8'h00;
14'h344a:data=8'h00;
14'h344b:data=8'h00;
14'h344c:data=8'h00;
14'h344d:data=8'h00;
14'h344e:data=8'h00;
14'h344f:data=8'h00;
14'h3450:data=8'h00;
14'h3451:data=8'h00;
14'h3452:data=8'h00;
14'h3453:data=8'h00;
14'h3454:data=8'h00;
14'h3455:data=8'h00;
14'h3456:data=8'h00;
14'h3457:data=8'h00;
14'h3458:data=8'h00;
14'h3459:data=8'h00;
14'h345a:data=8'h00;
14'h345b:data=8'h00;
14'h345c:data=8'h00;
14'h345d:data=8'h00;
14'h345e:data=8'h00;
14'h345f:data=8'h00;
14'h3460:data=8'h00;
14'h3461:data=8'h00;
14'h3462:data=8'h00;
14'h3463:data=8'h00;
14'h3464:data=8'h00;
14'h3465:data=8'h00;
14'h3466:data=8'h00;
14'h3467:data=8'h00;
14'h3468:data=8'h00;
14'h3469:data=8'h00;
14'h346a:data=8'h00;
14'h346b:data=8'h00;
14'h346c:data=8'h00;
14'h346d:data=8'h00;
14'h346e:data=8'h00;
14'h346f:data=8'h00;
14'h3470:data=8'h00;
14'h3471:data=8'h00;
14'h3472:data=8'h00;
14'h3473:data=8'h00;
14'h3474:data=8'h00;
14'h3475:data=8'h00;
14'h3476:data=8'h00;
14'h3477:data=8'h00;
14'h3478:data=8'h00;
14'h3479:data=8'h00;
14'h347a:data=8'h00;
14'h347b:data=8'h00;
14'h347c:data=8'h00;
14'h347d:data=8'h00;
14'h347e:data=8'h00;
14'h347f:data=8'h00;
14'h3c00:data=8'h00;
14'h3c01:data=8'h00;
14'h3c02:data=8'h00;
14'h3c03:data=8'h00;
14'h3c04:data=8'h00;
14'h3c05:data=8'h00;
14'h3c06:data=8'h00;
14'h3c07:data=8'h00;
14'h3c08:data=8'h00;
14'h3c09:data=8'h00;
14'h3c0a:data=8'h00;
14'h3c0b:data=8'h00;
14'h3c0c:data=8'h00;
14'h3c0d:data=8'h00;
14'h3c0e:data=8'h00;
14'h3c0f:data=8'h00;
14'h3c10:data=8'h00;
14'h3c11:data=8'h00;
14'h3c12:data=8'h00;
14'h3c13:data=8'h00;
14'h3c14:data=8'h00;
14'h3c15:data=8'h00;
14'h3c16:data=8'h00;
14'h3c17:data=8'h00;
14'h3c18:data=8'h00;
14'h3c19:data=8'h00;
14'h3c1a:data=8'h00;
14'h3c1b:data=8'h00;
14'h3c1c:data=8'h00;
14'h3c1d:data=8'h00;
14'h3c1e:data=8'h00;
14'h3c1f:data=8'h00;
14'h3c20:data=8'h00;
14'h3c21:data=8'h00;
14'h3c22:data=8'h00;
14'h3c23:data=8'h00;
14'h3c24:data=8'h00;
14'h3c25:data=8'h00;
14'h3c26:data=8'h00;
14'h3c27:data=8'h00;
14'h3c28:data=8'h00;
14'h3c29:data=8'h00;
14'h3c2a:data=8'h00;
14'h3c2b:data=8'h00;
14'h3c2c:data=8'h00;
14'h3c2d:data=8'h00;
14'h3c2e:data=8'h00;
14'h3c2f:data=8'h00;
14'h3c30:data=8'h00;
14'h3c31:data=8'h00;
14'h3c32:data=8'h00;
14'h3c33:data=8'h00;
14'h3c34:data=8'h00;
14'h3c35:data=8'h00;
14'h3c36:data=8'h00;
14'h3c37:data=8'h00;
14'h3c38:data=8'h00;
14'h3c39:data=8'h00;
14'h3c3a:data=8'h00;
14'h3c3b:data=8'h00;
14'h3c3c:data=8'h00;
14'h3c3d:data=8'h00;
14'h3c3e:data=8'h00;
14'h3c3f:data=8'h00;
14'h3c40:data=8'h00;
14'h3c41:data=8'h00;
14'h3c42:data=8'h00;
14'h3c43:data=8'h00;
14'h3c44:data=8'h00;
14'h3c45:data=8'h00;
14'h3c46:data=8'h00;
14'h3c47:data=8'h00;
14'h3c48:data=8'h00;
14'h3c49:data=8'h00;
14'h3c4a:data=8'h00;
14'h3c4b:data=8'h00;
14'h3c4c:data=8'h00;
14'h3c4d:data=8'h00;
14'h3c4e:data=8'h00;
14'h3c4f:data=8'h00;
14'h3c50:data=8'h00;
14'h3c51:data=8'h00;
14'h3c52:data=8'h00;
14'h3c53:data=8'h00;
14'h3c54:data=8'h00;
14'h3c55:data=8'h00;
14'h3c56:data=8'h00;
14'h3c57:data=8'h00;
14'h3c58:data=8'h00;
14'h3c59:data=8'h00;
14'h3c5a:data=8'h00;
14'h3c5b:data=8'h00;
14'h3c5c:data=8'h00;
14'h3c5d:data=8'h00;
14'h3c5e:data=8'h00;
14'h3c5f:data=8'h00;
14'h3c60:data=8'h00;
14'h3c61:data=8'h00;
14'h3c62:data=8'h00;
14'h3c63:data=8'h00;
14'h3c64:data=8'h00;
14'h3c65:data=8'h00;
14'h3c66:data=8'h00;
14'h3c67:data=8'h00;
14'h3c68:data=8'h00;
14'h3c69:data=8'h00;
14'h3c6a:data=8'h00;
14'h3c6b:data=8'h00;
14'h3c6c:data=8'h00;
14'h3c6d:data=8'h00;
14'h3c6e:data=8'h00;
14'h3c6f:data=8'h00;
14'h3c70:data=8'h00;
14'h3c71:data=8'h00;
14'h3c72:data=8'h00;
14'h3c73:data=8'h00;
14'h3c74:data=8'h00;
14'h3c75:data=8'h00;
14'h3c76:data=8'h00;
14'h3c77:data=8'h00;
14'h3c78:data=8'h00;
14'h3c79:data=8'h00;
14'h3c7a:data=8'h00;
14'h3c7b:data=8'h00;
14'h3c7c:data=8'h00;
14'h3c7d:data=8'h00;
14'h3c7e:data=8'h00;
14'h3c7f:data=8'h00;





		default:data=8'h00;
		endcase
	end
endmodule
